module KERNAL(
       input clk,
       input[11:0] addr,
       output reg[31:0] out
);

always@(posedge clk)
case(addr[10:0])
11'd0: out <= 32'b00000000000000000000000000000000;
11'd1: out <= 32'b00000000010100000000001010100101;
11'd2: out <= 32'b00000000010100000000000001000011;
11'd3: out <= 32'b00000000010100000000000001001101;
11'd4: out <= 32'b00000001111100000000000000000000;
11'd5: out <= 32'b00000000010100000000000001101110;
11'd6: out <= 32'b00000000010100000000000001110101;
11'd7: out <= 32'b00000001111100000000000000000000;
11'd8: out <= 32'b00000000010100000000000001111100;
11'd9: out <= 32'b00000000000000000000000000000000;
11'd10: out <= 32'b00000000000100000000000000000000;
11'd11: out <= 32'b00000000000101000000000000000000;
11'd12: out <= 32'b00000000000110000000000000000000;
11'd13: out <= 32'b00000000000111000000000000000000;
11'd14: out <= 32'b00000001111100000000000000000000;
11'd15: out <= 32'b00000000000000000000000000000000;
11'd16: out <= 32'b00000000011100000001111111110000;
11'd17: out <= 32'b00000000011000000000000000000000;
11'd18: out <= 32'b00000000011100000001111111110001;
11'd19: out <= 32'b00000000011001000000000000000000;
11'd20: out <= 32'b00000000011100000001111111110010;
11'd21: out <= 32'b00000000011010000000000000000000;
11'd22: out <= 32'b00000000011100000001111111110011;
11'd23: out <= 32'b00000000011011000000000000000000;
11'd24: out <= 32'b00000001111100000000000000000000;
11'd25: out <= 32'b00000000000000000000000000000000;
11'd26: out <= 32'b00000000011100000001111111110000;
11'd27: out <= 32'b00000000011000000000000000000000;
11'd28: out <= 32'b00000000011100000001111111110001;
11'd29: out <= 32'b00000000011001000000000000000000;
11'd30: out <= 32'b00000000011100000001111111110010;
11'd31: out <= 32'b00000000011010000000000000000000;
11'd32: out <= 32'b00000000011100000001111111110011;
11'd33: out <= 32'b00000000011011000000000000000000;
11'd34: out <= 32'b00000001111000000000000000001001;
11'd35: out <= 32'b00000001111100000000000000000000;
11'd36: out <= 32'b00000000000000000000000000000000;
11'd37: out <= 32'b00000000011100000001111111110100;
11'd38: out <= 32'b00000000011000000000000000000000;
11'd39: out <= 32'b00000000011100000001111111110101;
11'd40: out <= 32'b00000000011001000000000000000000;
11'd41: out <= 32'b00000000011100000001111111110110;
11'd42: out <= 32'b00000000011010000000000000000000;
11'd43: out <= 32'b00000000011100000001111111110111;
11'd44: out <= 32'b00000000011011000000000000000000;
11'd45: out <= 32'b00000001111000000000000000001001;
11'd46: out <= 32'b00000001111100000000000000000000;
11'd47: out <= 32'b00000000000000000000000000000000;
11'd48: out <= 32'b00000000011100000001111111110000;
11'd49: out <= 32'b00000001100000000000000000000000;
11'd50: out <= 32'b00000000011100000001111111110001;
11'd51: out <= 32'b00000001100001000000000000000000;
11'd52: out <= 32'b00000000011100000001111111110010;
11'd53: out <= 32'b00000001100010000000000000000000;
11'd54: out <= 32'b00000000011100000001111111110011;
11'd55: out <= 32'b00000001100011000000000000000000;
11'd56: out <= 32'b00000001111100000000000000000000;
11'd57: out <= 32'b00000000000000000000000000000000;
11'd58: out <= 32'b00000000011100000001111111110100;
11'd59: out <= 32'b00000001100000000000000000000000;
11'd60: out <= 32'b00000000011100000001111111110101;
11'd61: out <= 32'b00000001100001000000000000000000;
11'd62: out <= 32'b00000000011100000001111111110110;
11'd63: out <= 32'b00000001100010000000000000000000;
11'd64: out <= 32'b00000000011100000001111111110111;
11'd65: out <= 32'b00000001100011000000000000000000;
11'd66: out <= 32'b00000001111100000000000000000000;
11'd67: out <= 32'b00000000000000000000000000000000;
11'd68: out <= 32'b00000001111000000000000000100100;
11'd69: out <= 32'b00000000000011000000000000000010;
11'd70: out <= 32'b00000000001000000000000000000000;
11'd71: out <= 32'b00000000000101000000000000001111;
11'd72: out <= 32'b00000000110100010000000000000000;
11'd73: out <= 32'b00000000011100000001111111100000;
11'd74: out <= 32'b00000000011000000000000000000000;
11'd75: out <= 32'b00000001111000000000000000111001;
11'd76: out <= 32'b00000001111100000000000000000000;
11'd77: out <= 32'b00000000000000000000000000000000;
11'd78: out <= 32'b00000001111000000000000000100100;
11'd79: out <= 32'b00000000000011000000000000000011;
11'd80: out <= 32'b00000000001000000000000000000000;
11'd81: out <= 32'b00000000000101000000000011111111;
11'd82: out <= 32'b00000000110100010000000000000000;
11'd83: out <= 32'b00000000011100000001111111100001;
11'd84: out <= 32'b00000000011000000000000000000000;
11'd85: out <= 32'b00000001111000000000000000111001;
11'd86: out <= 32'b00000001111100000000000000000000;
11'd87: out <= 32'b00000000000000000000000000000000;
11'd88: out <= 32'b00000000000110000000000000000000;
11'd89: out <= 32'b00000000000111000001111111010000;
11'd90: out <= 32'b00000000000000000000000000000000;
11'd91: out <= 32'b00000000000100000000000000000011;
11'd92: out <= 32'b00000001100101100000000000000000;
11'd93: out <= 32'b00000001111000000000000010010100;
11'd94: out <= 32'b00000000000100000000000000000100;
11'd95: out <= 32'b00000000100111000000000000000000;
11'd96: out <= 32'b00000001100001000000000000000000;
11'd97: out <= 32'b00000001111000000000000010010100;
11'd98: out <= 32'b00000000000100001111111111100000;
11'd99: out <= 32'b00000000110101000000000000000000;
11'd100: out <= 32'b00000000000100000000000000000101;
11'd101: out <= 32'b00000001111000000000000010010100;
11'd102: out <= 32'b00000000010011000000000000000000;
11'd103: out <= 32'b00000000010010000000000000000000;
11'd104: out <= 32'b00000000000100000000000000000010;
11'd105: out <= 32'b00000001011110000000000000000000;
11'd106: out <= 32'b00000001010000000000000011100100;
11'd107: out <= 32'b00000000010100000000000011010111;
11'd108: out <= 32'b00000000000000000000000000000000;
11'd109: out <= 32'b00000001111100000000000000000000;
11'd110: out <= 32'b00000000000000000000000000000000;
11'd111: out <= 32'b00000001111000000000000000100100;
11'd112: out <= 32'b00000000011100000001111111000010;
11'd113: out <= 32'b00000000000100001111111111111111;
11'd114: out <= 32'b00000000011000000000000000000000;
11'd115: out <= 32'b00000001111000000000000000111001;
11'd116: out <= 32'b00000001111100000000000000000000;
11'd117: out <= 32'b00000000000000000000000000000000;
11'd118: out <= 32'b00000001111000000000000000100100;
11'd119: out <= 32'b00000000011100000001000000000010;
11'd120: out <= 32'b00000000000100001111111111111111;
11'd121: out <= 32'b00000000011000000000000000000000;
11'd122: out <= 32'b00000001111000000000000000111001;
11'd123: out <= 32'b00000001111100000000000000000000;
11'd124: out <= 32'b00000000000000000000000000000000;
11'd125: out <= 32'b00000001111100000000000000000000;
11'd126: out <= 32'b00000000000000000000000000000000;
11'd127: out <= 32'b00000001111000000000000000011001;
11'd128: out <= 32'b00000000000110000000000000000000;
11'd129: out <= 32'b00000000001110000000000000000000;
11'd130: out <= 32'b00000001111000000000000000101111;
11'd131: out <= 32'b00000001111100000000000000000000;
11'd132: out <= 32'b00000000000000000000000000000000;
11'd133: out <= 32'b00000001111000000000000000001111;
11'd134: out <= 32'b00000000000110000100000000000000;
11'd135: out <= 32'b00000000111000100000000000000000;
11'd136: out <= 32'b00000000001101000000000000000000;
11'd137: out <= 32'b00000000001100000000000000000001;
11'd138: out <= 32'b00000001111000000000000000101111;
11'd139: out <= 32'b00000001111100000000000000000000;
11'd140: out <= 32'b00000000000000000000000000000000;
11'd141: out <= 32'b00000001111000000000000000001111;
11'd142: out <= 32'b00000000000110001111000000000000;
11'd143: out <= 32'b00000000111000100000000000000000;
11'd144: out <= 32'b00000000001101000000000000000000;
11'd145: out <= 32'b00000000001100000000000000000001;
11'd146: out <= 32'b00000001111000000000000000101111;
11'd147: out <= 32'b00000001111100000000000000000000;
11'd148: out <= 32'b00000000000000000000000000000000;
11'd149: out <= 32'b00000001111000000000000000001111;
11'd150: out <= 32'b00000000000110001000000000000000;
11'd151: out <= 32'b00000000111000100000000000000000;
11'd152: out <= 32'b00000000001101000000000000000000;
11'd153: out <= 32'b00000000001100000000000000000001;
11'd154: out <= 32'b00000001111000000000000000101111;
11'd155: out <= 32'b00000001111100000000000000000000;
11'd156: out <= 32'b00000000000000000000000000000000;
11'd157: out <= 32'b00000000000100000001000000000000;
11'd158: out <= 32'b00000000000000000000000000000000;
11'd159: out <= 32'b00000000100100000000000000000000;
11'd160: out <= 32'b00000000000101000000000000000000;
11'd161: out <= 32'b00000000011001000000000000000000;
11'd162: out <= 32'b00000000010000000000000000000000;
11'd163: out <= 32'b00000000000101000010000000000000;
11'd164: out <= 32'b00000001011100010000000000000000;
11'd165: out <= 32'b00000001001000000000000010100111;
11'd166: out <= 32'b00000000010100000000000010011110;
11'd167: out <= 32'b00000000000000000000000000000000;
11'd168: out <= 32'b00000000000100000000000000000000;
11'd169: out <= 32'b00000000000101000000000000000000;
11'd170: out <= 32'b00000001111100000000000000000000;
11'd171: out <= 32'b00000000000000000000000000000000;
11'd172: out <= 32'b00000000000111000000111000000000;
11'd173: out <= 32'b00000000011100000001000000100000;
11'd174: out <= 32'b00000000000101000000000000000000;
11'd175: out <= 32'b00000000011001000000000000000000;
11'd176: out <= 32'b00000000000000000000000000000000;
11'd177: out <= 32'b00000000011100000001000000100000;
11'd178: out <= 32'b00000001100001000000000000000000;
11'd179: out <= 32'b00000000000100000000000000000110;
11'd180: out <= 32'b00000001111000000000000010010100;
11'd181: out <= 32'b00000000000110000000000000000000;
11'd182: out <= 32'b00000000000000000000000000000000;
11'd183: out <= 32'b00000000000100000000000000000111;
11'd184: out <= 32'b00000001100101100000000000000000;
11'd185: out <= 32'b00000001111000000000000010010100;
11'd186: out <= 32'b00000000100111000000000000000000;
11'd187: out <= 32'b00000001100001000000000000000000;
11'd188: out <= 32'b00000000000100000000000000001000;
11'd189: out <= 32'b00000001111000000000000010010100;
11'd190: out <= 32'b00000000000100000000000000001001;
11'd191: out <= 32'b00000001111000000000000010010100;
11'd192: out <= 32'b00000000010011000000000000000000;
11'd193: out <= 32'b00000000010010000000000000000000;
11'd194: out <= 32'b00000000000100000000000000000111;
11'd195: out <= 32'b00000001011110000000000000000000;
11'd196: out <= 32'b00000001010000000000000011000110;
11'd197: out <= 32'b00000000010100000000000010110110;
11'd198: out <= 32'b00000000000000000000000000000000;
11'd199: out <= 32'b00000000011100000001000000100000;
11'd200: out <= 32'b00000001100001000000000000000000;
11'd201: out <= 32'b00000000000100000000000000111111;
11'd202: out <= 32'b00000001011101000000000000000000;
11'd203: out <= 32'b00000001010000000000000011001111;
11'd204: out <= 32'b00000000010001000000000000000000;
11'd205: out <= 32'b00000000011001000000000000000000;
11'd206: out <= 32'b00000000010100000000000010110000;
11'd207: out <= 32'b00000000000000000000000000000000;
11'd208: out <= 32'b00000000011100000001000000100000;
11'd209: out <= 32'b00000000000100000000000000000000;
11'd210: out <= 32'b00000000011000000000000000000000;
11'd211: out <= 32'b00000001111000000000000000001001;
11'd212: out <= 32'b00000001111100000000000000000000;
11'd213: out <= 32'b00000000000000000000000000000000;
11'd214: out <= 32'b00000000000110000000000000000000;
11'd215: out <= 32'b00000000000000000000000000000000;
11'd216: out <= 32'b00000000000100000000000000000011;
11'd217: out <= 32'b00000001100101100000000000000000;
11'd218: out <= 32'b00000001111000000000000010010100;
11'd219: out <= 32'b00000000000100000000000000000100;
11'd220: out <= 32'b00000000000101000000000000000000;
11'd221: out <= 32'b00000001111000000000000010010100;
11'd222: out <= 32'b00000000010011000000000000000000;
11'd223: out <= 32'b00000000010010000000000000000000;
11'd224: out <= 32'b00000000000100000000000000000010;
11'd225: out <= 32'b00000001011110000000000000000000;
11'd226: out <= 32'b00000001010000000000000011100100;
11'd227: out <= 32'b00000000010100000000000011010111;
11'd228: out <= 32'b00000000000000000000000000000000;
11'd229: out <= 32'b00000001111100000000000000000000;
11'd230: out <= 32'b00000000000000000000000000000000;
11'd231: out <= 32'b00000000000000000000000000000000;
11'd232: out <= 32'b00000000011100000001000000000010;
11'd233: out <= 32'b00000001100000000000000000000000;
11'd234: out <= 32'b00000000000101001111111111111111;
11'd235: out <= 32'b00000001011100010000000000000000;
11'd236: out <= 32'b00000001001000000000000011101110;
11'd237: out <= 32'b00000000010100000000000011100111;
11'd238: out <= 32'b00000000000000000000000000000000;
11'd239: out <= 32'b00000001111100000000000000000000;
11'd240: out <= 32'b00000000000000000000000000000000;
11'd241: out <= 32'b00000001111000000000000000001001;
11'd242: out <= 32'b00000000011100000001000000000010;
11'd243: out <= 32'b00000000000100000000000000000000;
11'd244: out <= 32'b00000000011000000000000000000000;
11'd245: out <= 32'b00000000000100000000000011111101;
11'd246: out <= 32'b00000000000101000000000000000000;
11'd247: out <= 32'b00000001111000000000000010010100;
11'd248: out <= 32'b00000001111000000000000011100110;
11'd249: out <= 32'b00000001111100000000000000000000;
11'd250: out <= 32'b00000000000000000000000000000000;
11'd251: out <= 32'b00000001111000000000000000001001;
11'd252: out <= 32'b00000000011100000001111110100101;
11'd253: out <= 32'b00000000000111000000000000000000;
11'd254: out <= 32'b00000000011011000000000000000000;
11'd255: out <= 32'b00000000000110000001111110101000;
11'd256: out <= 32'b00000000000000000000000000000000;
11'd257: out <= 32'b00000000100110000000000000000000;
11'd258: out <= 32'b00000000000111000000000000000000;
11'd259: out <= 32'b00000000011011000000000000000000;
11'd260: out <= 32'b00000000010010000000000000000000;
11'd261: out <= 32'b00000000000101000001111110101101;
11'd262: out <= 32'b00000001011110010000000000000000;
11'd263: out <= 32'b00000001010100000000000100000000;
11'd264: out <= 32'b00000000011100000001111110101101;
11'd265: out <= 32'b00000000000111000000000000001111;
11'd266: out <= 32'b00000000011011000000000000000000;
11'd267: out <= 32'b00000000000000000000000000000000;
11'd268: out <= 32'b00000000011100000001111110100100;
11'd269: out <= 32'b00000001100000000000000000000000;
11'd270: out <= 32'b00000001100110000000000000000000;
11'd271: out <= 32'b00000000000101001000000000000000;
11'd272: out <= 32'b00000000110100010000000000000000;
11'd273: out <= 32'b00000000000101000000000000000111;
11'd274: out <= 32'b00000001000000010000000000000000;
11'd275: out <= 32'b00000001001100000000000000000000;
11'd276: out <= 32'b00000000000101000000000000000110;
11'd277: out <= 32'b00000001000000010000000000000000;
11'd278: out <= 32'b00000001001100000000000000000000;
11'd279: out <= 32'b00000001100111000000000000000000;
11'd280: out <= 32'b00000000000101000000000000000000;
11'd281: out <= 32'b00000000111110010000000000000000;
11'd282: out <= 32'b00000001001110000000000000000000;
11'd283: out <= 32'b00000000000101001111111111111111;
11'd284: out <= 32'b00000000110110010000000000000000;
11'd285: out <= 32'b00000000011010000000000000000000;
11'd286: out <= 32'b00000000011100000001111110101110;
11'd287: out <= 32'b00000000000100000001111110101101;
11'd288: out <= 32'b00000000011000000000000000000000;
11'd289: out <= 32'b00000000000000000000000000000000;
11'd290: out <= 32'b00000000011100000001111110101110;
11'd291: out <= 32'b00000001100000000000000000000000;
11'd292: out <= 32'b00000001011000000000000000000000;
11'd293: out <= 32'b00000000011000000000000000000000;
11'd294: out <= 32'b00000000100100000000000000000000;
11'd295: out <= 32'b00000001100000000000000000000000;
11'd296: out <= 32'b00000000000101000000000000000101;
11'd297: out <= 32'b00000001011100010000000000000000;
11'd298: out <= 32'b00000001001000000000000100101101;
11'd299: out <= 32'b00000001010000000000000100101101;
11'd300: out <= 32'b00000000010100000000000100110000;
11'd301: out <= 32'b00000000000000000000000000000000;
11'd302: out <= 32'b00000000000101000000000000000011;
11'd303: out <= 32'b00000000101100010000000000000000;
11'd304: out <= 32'b00000000000000000000000000000000;
11'd305: out <= 32'b00000001100110000000000000000000;
11'd306: out <= 32'b00000000000101000000000000001000;
11'd307: out <= 32'b00000000110110010000000000000000;
11'd308: out <= 32'b00000000000101000000000000000010;
11'd309: out <= 32'b00000001000010010000000000000000;
11'd310: out <= 32'b00000001001110000000000000000000;
11'd311: out <= 32'b00000000000101000000000000000000;
11'd312: out <= 32'b00000000111100010000000000000000;
11'd313: out <= 32'b00000001001100000000000000000000;
11'd314: out <= 32'b00000000101100110000000000000000;
11'd315: out <= 32'b00000000000101000000000000001111;
11'd316: out <= 32'b00000000110100010000000000000000;
11'd317: out <= 32'b00000001100111100000000000000000;
11'd318: out <= 32'b00000000011000000000000000000000;
11'd319: out <= 32'b00000000011100000001111110101110;
11'd320: out <= 32'b00000001100000000000000000000000;
11'd321: out <= 32'b00000000000101000001111110101001;
11'd322: out <= 32'b00000001011100010000000000000000;
11'd323: out <= 32'b00000001010000000000000100100001;
11'd324: out <= 32'b00000000011100000001111110101000;
11'd325: out <= 32'b00000001100000000000000000000000;
11'd326: out <= 32'b00000000000101000000000000000101;
11'd327: out <= 32'b00000001011100010000000000000000;
11'd328: out <= 32'b00000001001000000000000101001011;
11'd329: out <= 32'b00000001010000000000000101001011;
11'd330: out <= 32'b00000000010100000000000101001110;
11'd331: out <= 32'b00000000000000000000000000000000;
11'd332: out <= 32'b00000000000101000000000000000011;
11'd333: out <= 32'b00000000101100010000000000000000;
11'd334: out <= 32'b00000000000000000000000000000000;
11'd335: out <= 32'b00000001100110000000000000000000;
11'd336: out <= 32'b00000000000101000000000000000000;
11'd337: out <= 32'b00000000111100010000000000000000;
11'd338: out <= 32'b00000001001100000000000000000000;
11'd339: out <= 32'b00000000101100110000000000000000;
11'd340: out <= 32'b00000000000101000000000000001111;
11'd341: out <= 32'b00000000110100010000000000000000;
11'd342: out <= 32'b00000000011000000000000000000000;
11'd343: out <= 32'b00000000011100000001111110100101;
11'd344: out <= 32'b00000001100000000000000000000000;
11'd345: out <= 32'b00000000000101000000000000001110;
11'd346: out <= 32'b00000001011100010000000000000000;
11'd347: out <= 32'b00000001010000000000000101011111;
11'd348: out <= 32'b00000000010000000000000000000000;
11'd349: out <= 32'b00000000011000000000000000000000;
11'd350: out <= 32'b00000000010100000000000100001011;
11'd351: out <= 32'b00000000000000000000000000000000;
11'd352: out <= 32'b00000000011100000001111110101000;
11'd353: out <= 32'b00000001100011000000000000000000;
11'd354: out <= 32'b00000000010011000000000000000000;
11'd355: out <= 32'b00000000011011000000000000000000;
11'd356: out <= 32'b00000000011100000001111110101001;
11'd357: out <= 32'b00000001100011000000000000000000;
11'd358: out <= 32'b00000000010011000000000000000000;
11'd359: out <= 32'b00000000011011000000000000000000;
11'd360: out <= 32'b00000000011100000001111110101010;
11'd361: out <= 32'b00000001100011000000000000000000;
11'd362: out <= 32'b00000000010011000000000000000000;
11'd363: out <= 32'b00000000011011000000000000000000;
11'd364: out <= 32'b00000000011100000001111110101011;
11'd365: out <= 32'b00000001100011000000000000000000;
11'd366: out <= 32'b00000000010011000000000000000000;
11'd367: out <= 32'b00000000011011000000000000000000;
11'd368: out <= 32'b00000000011100000001111110101100;
11'd369: out <= 32'b00000001100011000000000000000000;
11'd370: out <= 32'b00000000010011000000000000000000;
11'd371: out <= 32'b00000000011011000000000000000000;
11'd372: out <= 32'b00000001111100000000000000000000;
11'd373: out <= 32'b00000000000000000000000000000000;
11'd374: out <= 32'b00000000011100000001111110100100;
11'd375: out <= 32'b00000001100000000000000000000000;
11'd376: out <= 32'b00000000000101000000000000000000;
11'd377: out <= 32'b00000001011100010000000000000000;
11'd378: out <= 32'b00000001010100000000000101111100;
11'd379: out <= 32'b00000000010100000000000110000001;
11'd380: out <= 32'b00000000000000000000000000000000;
11'd381: out <= 32'b00000000011100000001111110110001;
11'd382: out <= 32'b00000000000101000000000000001011;
11'd383: out <= 32'b00000000011001000000000000000000;
11'd384: out <= 32'b00000000010100000000000110000110;
11'd385: out <= 32'b00000000000000000000000000000000;
11'd386: out <= 32'b00000000011100000001111110110001;
11'd387: out <= 32'b00000000000101000000000000000000;
11'd388: out <= 32'b00000000011001000000000000000000;
11'd389: out <= 32'b00000000010100000000000110000110;
11'd390: out <= 32'b00000000000000000000000000000000;
11'd391: out <= 32'b00000000011100000001111110100100;
11'd392: out <= 32'b00000001111000000000001001101011;
11'd393: out <= 32'b00000000011000000000000000000000;
11'd394: out <= 32'b00000001111000000000000011111010;
11'd395: out <= 32'b00000000011100000001111110101000;
11'd396: out <= 32'b00000001100000000000000000000000;
11'd397: out <= 32'b00000000011100000001111110110010;
11'd398: out <= 32'b00000000011000000000000000000000;
11'd399: out <= 32'b00000000011100000001111110101001;
11'd400: out <= 32'b00000001100000000000000000000000;
11'd401: out <= 32'b00000000011100000001111110110011;
11'd402: out <= 32'b00000000011000000000000000000000;
11'd403: out <= 32'b00000000011100000001111110101010;
11'd404: out <= 32'b00000001100000000000000000000000;
11'd405: out <= 32'b00000000011100000001111110110100;
11'd406: out <= 32'b00000000011000000000000000000000;
11'd407: out <= 32'b00000000011100000001111110101011;
11'd408: out <= 32'b00000001100000000000000000000000;
11'd409: out <= 32'b00000000011100000001111110110101;
11'd410: out <= 32'b00000000011000000000000000000000;
11'd411: out <= 32'b00000000011100000001111110101100;
11'd412: out <= 32'b00000001100000000000000000000000;
11'd413: out <= 32'b00000000011100000001111110110110;
11'd414: out <= 32'b00000000011000000000000000000000;
11'd415: out <= 32'b00000000011100000001111110110111;
11'd416: out <= 32'b00000000000100000000000000001111;
11'd417: out <= 32'b00000000011000000000000000000000;
11'd418: out <= 32'b00000001111000000000000111110011;
11'd419: out <= 32'b00000001111100000000000000000000;
11'd420: out <= 32'b00000000000000000000000000000000;
11'd421: out <= 32'b00000000011100000001111110110000;
11'd422: out <= 32'b00000001100000000000000000000000;
11'd423: out <= 32'b00000000000101000000000000000000;
11'd424: out <= 32'b00000001011100010000000000000000;
11'd425: out <= 32'b00000001010100000000000110101011;
11'd426: out <= 32'b00000000010100000000000110110000;
11'd427: out <= 32'b00000000000000000000000000000000;
11'd428: out <= 32'b00000000011100000001111110110001;
11'd429: out <= 32'b00000000000101000000000000001011;
11'd430: out <= 32'b00000000011001000000000000000000;
11'd431: out <= 32'b00000000010100000000000110110101;
11'd432: out <= 32'b00000000000000000000000000000000;
11'd433: out <= 32'b00000000011100000001111110110001;
11'd434: out <= 32'b00000000000101000000000000000000;
11'd435: out <= 32'b00000000011001000000000000000000;
11'd436: out <= 32'b00000000010100000000000110110101;
11'd437: out <= 32'b00000000000000000000000000000000;
11'd438: out <= 32'b00000000011100000001111110110000;
11'd439: out <= 32'b00000001111000000000001001101011;
11'd440: out <= 32'b00000000011000000000000000000000;
11'd441: out <= 32'b00000001100000000000000000000000;
11'd442: out <= 32'b00000000000101000000000011111111;
11'd443: out <= 32'b00000000110100010000000000000000;
11'd444: out <= 32'b00000000011100000001111110100100;
11'd445: out <= 32'b00000000000101000000000000000111;
11'd446: out <= 32'b00000000111100010000000000000000;
11'd447: out <= 32'b00000001001100000000000000000000;
11'd448: out <= 32'b00000000000101000010011100010000;
11'd449: out <= 32'b00000001110000010000000000000001;
11'd450: out <= 32'b00000001001100000000000000000000;
11'd451: out <= 32'b00000000011000000000000000000000;
11'd452: out <= 32'b00000001111000000000000011111010;
11'd453: out <= 32'b00000000011100000001111110110101;
11'd454: out <= 32'b00000000000100000000000000111010;
11'd455: out <= 32'b00000000011000000000000000000000;
11'd456: out <= 32'b00000000011100000001111110101001;
11'd457: out <= 32'b00000001100000000000000000000000;
11'd458: out <= 32'b00000000011100000001111110110110;
11'd459: out <= 32'b00000000011000000000000000000000;
11'd460: out <= 32'b00000000011100000001111110101010;
11'd461: out <= 32'b00000001100000000000000000000000;
11'd462: out <= 32'b00000000011100000001111110110111;
11'd463: out <= 32'b00000000011000000000000000000000;
11'd464: out <= 32'b00000000011100000001111110101011;
11'd465: out <= 32'b00000001100000000000000000000000;
11'd466: out <= 32'b00000000011100000001111110111000;
11'd467: out <= 32'b00000000011000000000000000000000;
11'd468: out <= 32'b00000000011100000001111110101100;
11'd469: out <= 32'b00000001100000000000000000000000;
11'd470: out <= 32'b00000000011100000001111110111001;
11'd471: out <= 32'b00000000011000000000000000000000;
11'd472: out <= 32'b00000000011100000001111110111010;
11'd473: out <= 32'b00000000000100000000000000001111;
11'd474: out <= 32'b00000000011000000000000000000000;
11'd475: out <= 32'b00000000011100000001111110110000;
11'd476: out <= 32'b00000001100000000000000000000000;
11'd477: out <= 32'b00000000000101001111111100000000;
11'd478: out <= 32'b00000000110100010000000000000000;
11'd479: out <= 32'b00000000000101000000000000000111;
11'd480: out <= 32'b00000001000000010000000000000000;
11'd481: out <= 32'b00000001001100000000000000000000;
11'd482: out <= 32'b00000000011100000001111110100100;
11'd483: out <= 32'b00000000011000000000000000000000;
11'd484: out <= 32'b00000001111000000000000011111010;
11'd485: out <= 32'b00000000011100000001111110101010;
11'd486: out <= 32'b00000001100000000000000000000000;
11'd487: out <= 32'b00000000011100000001111110110010;
11'd488: out <= 32'b00000000011000000000000000000000;
11'd489: out <= 32'b00000000011100000001111110101011;
11'd490: out <= 32'b00000001100000000000000000000000;
11'd491: out <= 32'b00000000011100000001111110110011;
11'd492: out <= 32'b00000000011000000000000000000000;
11'd493: out <= 32'b00000000011100000001111110101100;
11'd494: out <= 32'b00000001100000000000000000000000;
11'd495: out <= 32'b00000000011100000001111110110100;
11'd496: out <= 32'b00000000011000000000000000000000;
11'd497: out <= 32'b00000001111000000000000111110011;
11'd498: out <= 32'b00000001111100000000000000000000;
11'd499: out <= 32'b00000000000000000000000000000000;
11'd500: out <= 32'b00000000000000000000000000000000;
11'd501: out <= 32'b00000000011100000001111110110011;
11'd502: out <= 32'b00000001100000000000000000000000;
11'd503: out <= 32'b00000000000101000000000000111010;
11'd504: out <= 32'b00000001011100010000000000000000;
11'd505: out <= 32'b00000001001000000000001000101011;
11'd506: out <= 32'b00000000000101000000000000001111;
11'd507: out <= 32'b00000001011100010000000000000000;
11'd508: out <= 32'b00000001001000000000001000101011;
11'd509: out <= 32'b00000000011100000001111110110010;
11'd510: out <= 32'b00000001100000000000000000000000;
11'd511: out <= 32'b00000000000101000000000000000000;
11'd512: out <= 32'b00000001011100010000000000000000;
11'd513: out <= 32'b00000001001000000000001000000110;
11'd514: out <= 32'b00000000000101000000000000000001;
11'd515: out <= 32'b00000001011100010000000000000000;
11'd516: out <= 32'b00000001001000000000001000000110;
11'd517: out <= 32'b00000000010100000000001000101011;
11'd518: out <= 32'b00000000000000000000000000000000;
11'd519: out <= 32'b00000000011100000001111110110011;
11'd520: out <= 32'b00000001100011000000000000000000;
11'd521: out <= 32'b00000000011100000001111110110010;
11'd522: out <= 32'b00000000011011000000000000000000;
11'd523: out <= 32'b00000000011100000001111110110100;
11'd524: out <= 32'b00000001100011000000000000000000;
11'd525: out <= 32'b00000000011100000001111110110011;
11'd526: out <= 32'b00000000011011000000000000000000;
11'd527: out <= 32'b00000000011100000001111110110101;
11'd528: out <= 32'b00000001100011000000000000000000;
11'd529: out <= 32'b00000000011100000001111110110100;
11'd530: out <= 32'b00000000011011000000000000000000;
11'd531: out <= 32'b00000000011100000001111110110110;
11'd532: out <= 32'b00000001100011000000000000000000;
11'd533: out <= 32'b00000000011100000001111110110101;
11'd534: out <= 32'b00000000011011000000000000000000;
11'd535: out <= 32'b00000000011100000001111110110111;
11'd536: out <= 32'b00000001100011000000000000000000;
11'd537: out <= 32'b00000000011100000001111110110110;
11'd538: out <= 32'b00000000011011000000000000000000;
11'd539: out <= 32'b00000000011100000001111110111000;
11'd540: out <= 32'b00000001100011000000000000000000;
11'd541: out <= 32'b00000000011100000001111110110111;
11'd542: out <= 32'b00000000011011000000000000000000;
11'd543: out <= 32'b00000000011100000001111110111001;
11'd544: out <= 32'b00000001100011000000000000000000;
11'd545: out <= 32'b00000000011100000001111110111000;
11'd546: out <= 32'b00000000011011000000000000000000;
11'd547: out <= 32'b00000000011100000001111110111010;
11'd548: out <= 32'b00000001100011000000000000000000;
11'd549: out <= 32'b00000000011100000001111110111001;
11'd550: out <= 32'b00000000011011000000000000000000;
11'd551: out <= 32'b00000000011100000001111110111010;
11'd552: out <= 32'b00000000000111000000000000000000;
11'd553: out <= 32'b00000000011011000000000000000000;
11'd554: out <= 32'b00000000010100000000000111110100;
11'd555: out <= 32'b00000000000000000000000000000000;
11'd556: out <= 32'b00000001111100000000000000000000;
11'd557: out <= 32'b00000000000000000000000000000000;
11'd558: out <= 32'b00000001111000000000000000001001;
11'd559: out <= 32'b00000000000111000000000000000000;
11'd560: out <= 32'b00000000000000000000000000000000;
11'd561: out <= 32'b00000000000100000000000000001010;
11'd562: out <= 32'b00000000011100000001111111000000;
11'd563: out <= 32'b00000001100001000000000000000000;
11'd564: out <= 32'b00000000000110000000000000000010;
11'd565: out <= 32'b00000000111101100000000000000000;
11'd566: out <= 32'b00000001001101000000000000000000;
11'd567: out <= 32'b00000001111000000000000010010100;
11'd568: out <= 32'b00000000000100000000000000001011;
11'd569: out <= 32'b00000000011100000001111111000001;
11'd570: out <= 32'b00000001100001000000000000000000;
11'd571: out <= 32'b00000000000110000000000000000010;
11'd572: out <= 32'b00000000111101100000000000000000;
11'd573: out <= 32'b00000001001101000000000000000000;
11'd574: out <= 32'b00000001111000000000000010010100;
11'd575: out <= 32'b00000000000100000000000000001100;
11'd576: out <= 32'b00000000011100000001111111000011;
11'd577: out <= 32'b00000001100001000000000000000000;
11'd578: out <= 32'b00000001100110010000000000000000;
11'd579: out <= 32'b00000000010010000000000000000000;
11'd580: out <= 32'b00000000011010000000000000000000;
11'd581: out <= 32'b00000000100101000000000000000000;
11'd582: out <= 32'b00000001100001000000000000000000;
11'd583: out <= 32'b00000000000110000000000011111111;
11'd584: out <= 32'b00000000110101100000000000000000;
11'd585: out <= 32'b00000000000110000000000000011111;
11'd586: out <= 32'b00000001011101100000000000000000;
11'd587: out <= 32'b00000001001000000000001001010110;
11'd588: out <= 32'b00000000000110000000000000001111;
11'd589: out <= 32'b00000001011101100000000000000000;
11'd590: out <= 32'b00000001001000000000001001101001;
11'd591: out <= 32'b00000001111000000000000010010100;
11'd592: out <= 32'b00000000011100000001111111000000;
11'd593: out <= 32'b00000001100001000000000000000000;
11'd594: out <= 32'b00000000000110000000000000100000;
11'd595: out <= 32'b00000001011101100000000000000000;
11'd596: out <= 32'b00000001010000000000001001010110;
11'd597: out <= 32'b00000000010100000000001001011110;
11'd598: out <= 32'b00000000000000000000000000000000;
11'd599: out <= 32'b00000000011100000001111111000000;
11'd600: out <= 32'b00000000000101000000000000000100;
11'd601: out <= 32'b00000000011001000000000000000000;
11'd602: out <= 32'b00000000011100000001111111000001;
11'd603: out <= 32'b00000001100001000000000000000000;
11'd604: out <= 32'b00000000010001000000000000000000;
11'd605: out <= 32'b00000000011001000000000000000000;
11'd606: out <= 32'b00000000000000000000000000000000;
11'd607: out <= 32'b00000000011100000001111111000000;
11'd608: out <= 32'b00000001100001000000000000000000;
11'd609: out <= 32'b00000000010001000000000000000000;
11'd610: out <= 32'b00000000011001000000000000000000;
11'd611: out <= 32'b00000000010011000000000000000000;
11'd612: out <= 32'b00000000000101000000000000111010;
11'd613: out <= 32'b00000001011111010000000000000000;
11'd614: out <= 32'b00000001001000000000001001101001;
11'd615: out <= 32'b00000001010000000000001001101001;
11'd616: out <= 32'b00000000010100000000001000110000;
11'd617: out <= 32'b00000000000000000000000000000000;
11'd618: out <= 32'b00000001111100000000000000000000;
11'd619: out <= 32'b00000000000000000000000000000000;
11'd620: out <= 32'b00000000000101000000000000000000;
11'd621: out <= 32'b00000001011100010000000000000000;
11'd622: out <= 32'b00000001010100000000001001110000;
11'd623: out <= 32'b00000000010100000000001001110011;
11'd624: out <= 32'b00000000000000000000000000000000;
11'd625: out <= 32'b00000000101000000000000000000000;
11'd626: out <= 32'b00000000010000000000000000000000;
11'd627: out <= 32'b00000000000000000000000000000000;
11'd628: out <= 32'b00000001111100000000000000000000;
11'd629: out <= 32'b00000000000000000000000000000000;
11'd630: out <= 32'b00000001110000010000000000000000;
11'd631: out <= 32'b00000001001110000000000000000000;
11'd632: out <= 32'b00000001110000010000000000000001;
11'd633: out <= 32'b00000001001111000000000000000000;
11'd634: out <= 32'b00000000000100001111111100000000;
11'd635: out <= 32'b00000000110110000000000000000000;
11'd636: out <= 32'b00000000000100000000000011111111;
11'd637: out <= 32'b00000000110111000000000000000000;
11'd638: out <= 32'b00000000000100000000000000000111;
11'd639: out <= 32'b00000001000010000000000000000000;
11'd640: out <= 32'b00000001001110000000000000000000;
11'd641: out <= 32'b00000000111111000000000000000000;
11'd642: out <= 32'b00000001001111000000000000000000;
11'd643: out <= 32'b00000000111011100000000000000000;
11'd644: out <= 32'b00000001100100110000000000000000;
11'd645: out <= 32'b00000001111100000000000000000000;
11'd646: out <= 32'b00000000000000000000000000000000;
11'd647: out <= 32'b00000000000000000000000000000000;
11'd648: out <= 32'b00000000000110000000000011111111;
11'd649: out <= 32'b00000001011100100000000000000000;
11'd650: out <= 32'b00000001010000000000001010001110;
11'd651: out <= 32'b00000001011101100000000000000000;
11'd652: out <= 32'b00000001010000000000001010001110;
11'd653: out <= 32'b00000000010100000000001010010101;
11'd654: out <= 32'b00000000000000000000000000000000;
11'd655: out <= 32'b00000000000110000000000000000000;
11'd656: out <= 32'b00000001000000100000000000000000;
11'd657: out <= 32'b00000001001100000000000000000000;
11'd658: out <= 32'b00000001000001100000000000000000;
11'd659: out <= 32'b00000001001101000000000000000000;
11'd660: out <= 32'b00000000010100000000001010000111;
11'd661: out <= 32'b00000000000000000000000000000000;
11'd662: out <= 32'b00000001110100010000000000000000;
11'd663: out <= 32'b00000001001110000000000000000000;
11'd664: out <= 32'b00000001110100010000000000000001;
11'd665: out <= 32'b00000001001111000000000000000000;
11'd666: out <= 32'b00000000000100000000000000000111;
11'd667: out <= 32'b00000000111111000000000000000000;
11'd668: out <= 32'b00000001001111000000000000000000;
11'd669: out <= 32'b00000001110111010000000000000000;
11'd670: out <= 32'b00000001001111000000000000000000;
11'd671: out <= 32'b00000000000100000000000000000111;
11'd672: out <= 32'b00000000111110000000000000000000;
11'd673: out <= 32'b00000001001110000000000000000000;
11'd674: out <= 32'b00000001100100100000000000000000;
11'd675: out <= 32'b00000000111000110000000000000000;
11'd676: out <= 32'b00000001111100000000000000000000;
11'd677: out <= 32'b00000000000000000000000000000000;
11'd678: out <= 32'b00000001111000000000000010011100;
11'd679: out <= 32'b00000001111000000000000011010101;
11'd680: out <= 32'b00000001111000000000000010101011;
11'd681: out <= 32'b00000000000100000000001101000000;
11'd682: out <= 32'b00000000011100000001111111010000;
11'd683: out <= 32'b00000000011000000000000000000000;
11'd684: out <= 32'b00000000011100000001111110101111;
11'd685: out <= 32'b00000000000111000000000000000000;
11'd686: out <= 32'b00000000011011000000000000000000;
11'd687: out <= 32'b00000001111000000000000001010111;
11'd688: out <= 32'b00000001111000000000000000001001;
11'd689: out <= 32'b00000000010100000000001011010000;
11'd690: out <= 32'b00000000000000000000000000000000;
11'd691: out <= 32'b00000000011100000001000000010000;
11'd692: out <= 32'b00000001100000000000000000000000;
11'd693: out <= 32'b00000000000101000000000000001111;
11'd694: out <= 32'b00000001011100010000000000000000;
11'd695: out <= 32'b00000001001000000000001011001011;
11'd696: out <= 32'b00000001100101000000000000000000;
11'd697: out <= 32'b00000000010001000000000000000000;
11'd698: out <= 32'b00000000011100000001000000010000;
11'd699: out <= 32'b00000000011001000000000000000000;
11'd700: out <= 32'b00000000000110000000000000000111;
11'd701: out <= 32'b00000001011101100000000000000000;
11'd702: out <= 32'b00000001010100000000001011000000;
11'd703: out <= 32'b00000000010100000000001011000100;
11'd704: out <= 32'b00000000000000000000000000000000;
11'd705: out <= 32'b00000000000100000000000000000001;
11'd706: out <= 32'b00000000000101000000000000001111;
11'd707: out <= 32'b00000000010100000000001011001000;
11'd708: out <= 32'b00000000000000000000000000000000;
11'd709: out <= 32'b00000000000100000000000000000001;
11'd710: out <= 32'b00000000000101000000000000000010;
11'd711: out <= 32'b00000000010100000000001011001000;
11'd712: out <= 32'b00000000000000000000000000000000;
11'd713: out <= 32'b00000001111000000000000010001100;
11'd714: out <= 32'b00000001111100000000000000000000;
11'd715: out <= 32'b00000000000000000000000000000000;
11'd716: out <= 32'b00000000000100000000000000000010;
11'd717: out <= 32'b00000000000101000000000000000000;
11'd718: out <= 32'b00000001111000000000000010001100;
11'd719: out <= 32'b00000001111100000000000000000000;
11'd720: out <= 32'b00000000000000000000000000000000;
11'd721: out <= 32'b00000001111000000000000011110000;
11'd722: out <= 32'b00000000011100000001111111000000;
11'd723: out <= 32'b00000000000101000000000000000101;
11'd724: out <= 32'b00000000011001000000000000000000;
11'd725: out <= 32'b00000000011100000001111111000001;
11'd726: out <= 32'b00000000000101000000000000000011;
11'd727: out <= 32'b00000000011001000000000000000000;
11'd728: out <= 32'b00000000011100000001111111000011;
11'd729: out <= 32'b00000000000101000000110100000000;
11'd730: out <= 32'b00000000011001000000000000000000;
11'd731: out <= 32'b00000001111000000000001000101101;
11'd732: out <= 32'b00000000000100001111111111111111;
11'd733: out <= 32'b00000000011100000001111110110000;
11'd734: out <= 32'b00000000011000000000000000000000;
11'd735: out <= 32'b00000001111000000000000110100100;
11'd736: out <= 32'b00000000011100000001111111000011;
11'd737: out <= 32'b00000000000101000001111110110001;
11'd738: out <= 32'b00000000011001000000000000000000;
11'd739: out <= 32'b00000001111000000000001000101101;
11'd740: out <= 32'b00000000011100000001111111000001;
11'd741: out <= 32'b00000000000101000000000000000100;
11'd742: out <= 32'b00000000011001000000000000000000;
11'd743: out <= 32'b00000000011100000001111111100001;
11'd744: out <= 32'b00000001100000000000000000000000;
11'd745: out <= 32'b00000000011100000001111110100100;
11'd746: out <= 32'b00000000011000000000000000000000;
11'd747: out <= 32'b00000000011100000001111111100001;
11'd748: out <= 32'b00000000000101000000000000000000;
11'd749: out <= 32'b00000000011000000000000000000000;
11'd750: out <= 32'b00000001111000000000000101110101;
11'd751: out <= 32'b00000000011100000001111111000000;
11'd752: out <= 32'b00000001100001000000000000000000;
11'd753: out <= 32'b00000000010001000000000000000000;
11'd754: out <= 32'b00000000011001000000000000000000;
11'd755: out <= 32'b00000000011100000001111111000011;
11'd756: out <= 32'b00000000000101000001111110110001;
11'd757: out <= 32'b00000000011001000000000000000000;
11'd758: out <= 32'b00000001111000000000001000101101;
11'd759: out <= 32'b00000001111000000000000000001001;
11'd760: out <= 32'b00000000000100000000000000001101;
11'd761: out <= 32'b00000000000101000000000000000001;
11'd762: out <= 32'b00000001111000000000000010010100;
11'd763: out <= 32'b00000001111000000000001010110010;
11'd764: out <= 32'b00000000000100000000000000000101;
11'd765: out <= 32'b00000000000101000000000000000000;
11'd766: out <= 32'b00000001111000000000000010000100;
11'd767: out <= 32'b00000000011100000001111111000010;
11'd768: out <= 32'b00000000000100000000000000000000;
11'd769: out <= 32'b00000000011000000000000000000000;
11'd770: out <= 32'b00000000000000000000000000000000;
11'd771: out <= 32'b00000001100000000000000000000000;
11'd772: out <= 32'b00000000000101001111111111111111;
11'd773: out <= 32'b00000001011100010000000000000000;
11'd774: out <= 32'b00000001001000000000001100001000;
11'd775: out <= 32'b00000000010100000000001100000010;
11'd776: out <= 32'b00000000000000000000000000000000;
11'd777: out <= 32'b00000000000101000000000000000000;
11'd778: out <= 32'b00000000011001000000000000000000;
11'd779: out <= 32'b00000000010100000000001011010000;
11'd780: out <= 32'b11010101101111111010101000010101;
11'd781: out <= 32'b11111010110101000010111000011000;
11'd782: out <= 32'b01101100100101100000110000000101;
11'd783: out <= 32'b01111110000111000111001000001101;
11'd784: out <= 32'b01100110000011011011110111101010;
11'd785: out <= 32'b10101100100101000100011100010000;
11'd786: out <= 32'b10011101000101001111111111111010;
11'd787: out <= 32'b00000011001001001101110100100011;
11'd788: out <= 32'b10111110100010110100110010110111;
11'd789: out <= 32'b10111000101010011100001101000100;
11'd790: out <= 32'b11100101001000000010011001011101;
11'd791: out <= 32'b10000110100000110001110101101011;
11'd792: out <= 32'b10101100110011000000011111010110;
11'd793: out <= 32'b01000011110010000010001100111000;
11'd794: out <= 32'b00101001101110101100110101101110;
11'd795: out <= 32'b11110101000001011001110110010110;
11'd796: out <= 32'b11111011101011110010011000001001;
11'd797: out <= 32'b01001010110010100000000010011011;
11'd798: out <= 32'b10010111110110010001100010010011;
11'd799: out <= 32'b01101101000101101011011000110100;
11'd800: out <= 32'b11110100001110011011100101001101;
11'd801: out <= 32'b00110000101000101110100101000000;
11'd802: out <= 32'b00110000100110100110101000011100;
11'd803: out <= 32'b01111110110100111010111101000110;
11'd804: out <= 32'b01011000101010110011010011011101;
11'd805: out <= 32'b11110001001110100111001000011010;
11'd806: out <= 32'b00010011010000000110110011101011;
11'd807: out <= 32'b01001001011101111101110110101100;
11'd808: out <= 32'b00100010111111100110101101001000;
11'd809: out <= 32'b00011000010011001100111101010011;
11'd810: out <= 32'b01111110110011011101111011101000;
11'd811: out <= 32'b11010100101011001010110100111000;
11'd812: out <= 32'b11100101010100110000110000000111;
11'd813: out <= 32'b10000001101110001110000110111100;
11'd814: out <= 32'b11100011101000010011111100011111;
11'd815: out <= 32'b11110011011111010100111011010100;
11'd816: out <= 32'b01101110000010101101001011111101;
11'd817: out <= 32'b01101101101001100110010011111111;
11'd818: out <= 32'b01100110001101100010101110000100;
11'd819: out <= 32'b01000011111101000110000100001011;
11'd820: out <= 32'b10001111000100010001010000000010;
11'd821: out <= 32'b11000110101111000001001011000010;
11'd822: out <= 32'b00100010111110000011100011000111;
11'd823: out <= 32'b00001010001010111011001111001101;
11'd824: out <= 32'b11001001000100100000100000101000;
11'd825: out <= 32'b11111100111010110000001000110110;
11'd826: out <= 32'b10000000110010000101100111101111;
11'd827: out <= 32'b11010110011011001111000001011111;
11'd828: out <= 32'b11011101101110101101010011011100;
11'd829: out <= 32'b00111010011100011010101001001110;
11'd830: out <= 32'b10011010110100110111111011100000;
11'd831: out <= 32'b01101111111101000111101111100000;
11'd832: out <= 32'b01100100001001100111100111111100;
11'd833: out <= 32'b01111000011101110100100011111101;
11'd834: out <= 32'b01100101100111101111001110010000;
11'd835: out <= 32'b11011000101001000110111111010011;
11'd836: out <= 32'b01001110110111100001010101000101;
11'd837: out <= 32'b01001011010110011110010011010101;
11'd838: out <= 32'b10101100110111111110101100100010;
11'd839: out <= 32'b10110011110001101000011111000000;
11'd840: out <= 32'b11001111001101011100010011001001;
11'd841: out <= 32'b01010101101001110001001000011101;
11'd842: out <= 32'b01010011001100111001110111100101;
11'd843: out <= 32'b10010101100101001010111000000010;
11'd844: out <= 32'b10111101011000000110100100101101;
11'd845: out <= 32'b00000100110000111001010110101100;
11'd846: out <= 32'b10001001101100010110100101000001;
11'd847: out <= 32'b11000000110011100011010100001101;
11'd848: out <= 32'b10111000010010100100000110011001;
11'd849: out <= 32'b01010110011010110011000100110011;
11'd850: out <= 32'b11101101001010000101000101100000;
11'd851: out <= 32'b10101011100101010100100001100100;
11'd852: out <= 32'b00000101111111101110110111011100;
11'd853: out <= 32'b01011110011100100101100010001111;
11'd854: out <= 32'b01101101111010100100000000011000;
11'd855: out <= 32'b10000110111111010100000100110100;
11'd856: out <= 32'b00010010110111001100010011000011;
11'd857: out <= 32'b10000101110001101101101010111100;
11'd858: out <= 32'b10101000001011000111110011100010;
11'd859: out <= 32'b11010011110010010110110111100111;
11'd860: out <= 32'b10000001001010110111000010100011;
11'd861: out <= 32'b11110000111100110000000001011001;
11'd862: out <= 32'b00111000000010010011010011000101;
11'd863: out <= 32'b10000110000000000010101101111101;
11'd864: out <= 32'b10001011100010000110011010010101;
11'd865: out <= 32'b00011011000110011110101010001011;
11'd866: out <= 32'b01011101010100010101110100110111;
11'd867: out <= 32'b11101111000010100001100011000000;
11'd868: out <= 32'b11011110000010011000011010011101;
11'd869: out <= 32'b10000100000010011000010001000100;
11'd870: out <= 32'b10011111110111011001101001001011;
11'd871: out <= 32'b00100001110110111100101111100011;
11'd872: out <= 32'b11011100101011001011101110100101;
11'd873: out <= 32'b10111010001111101100110011001100;
11'd874: out <= 32'b00010101111010011101000101000110;
11'd875: out <= 32'b01101001001010001001001101111001;
11'd876: out <= 32'b00010010100000100101011111101100;
11'd877: out <= 32'b01110001110001001011111000000100;
11'd878: out <= 32'b01111011100101000001001111110110;
11'd879: out <= 32'b01011000100001100010000101100011;
11'd880: out <= 32'b11110001000001010100100100001011;
11'd881: out <= 32'b00000110100101110111000000010101;
11'd882: out <= 32'b01111011101101111011110111001111;
11'd883: out <= 32'b00110110101101001111111110111000;
11'd884: out <= 32'b01001111001001110010000011011101;
11'd885: out <= 32'b11001100110111101100101011100000;
11'd886: out <= 32'b11000101101000111011011101001111;
11'd887: out <= 32'b10101110101000110101000010101100;
11'd888: out <= 32'b00101110000011011100010011000011;
11'd889: out <= 32'b10100111111000010101011110000011;
11'd890: out <= 32'b01011111001110000110010001010001;
11'd891: out <= 32'b01100000111010001100000101010011;
11'd892: out <= 32'b00101001010001010110111100000100;
11'd893: out <= 32'b11110101110001111001000001101001;
11'd894: out <= 32'b00101011110101110111111111011110;
11'd895: out <= 32'b11101011000001011110110100111011;
11'd896: out <= 32'b00100111100111011111000101101100;
11'd897: out <= 32'b00101100100010000011001010011100;
11'd898: out <= 32'b01001100001101010011101001010110;
11'd899: out <= 32'b01011000010100001111000011110010;
11'd900: out <= 32'b11011000101100001100010111101010;
11'd901: out <= 32'b01110101011001111100001010011010;
11'd902: out <= 32'b01011000001111000010111011011101;
11'd903: out <= 32'b11110001011010010101011101001010;
11'd904: out <= 32'b11011011000011001111010001001111;
11'd905: out <= 32'b01010011001000101110000001100101;
11'd906: out <= 32'b01101001110000011000001010101110;
11'd907: out <= 32'b10001000000110011100000100001011;
11'd908: out <= 32'b00000010001110001001110000000011;
11'd909: out <= 32'b01101101011000001010111010001110;
11'd910: out <= 32'b10101010010000010111110011000001;
11'd911: out <= 32'b10110001011010101101001011001001;
11'd912: out <= 32'b01110111110100000001111011101110;
11'd913: out <= 32'b01001001101100100111111010001100;
11'd914: out <= 32'b11111010101011110110110010011010;
11'd915: out <= 32'b00101110110001101110101000011111;
11'd916: out <= 32'b11001100001011001000000111101011;
11'd917: out <= 32'b11001010011001000000100000111011;
11'd918: out <= 32'b00001001101011011001000100010100;
11'd919: out <= 32'b11111111111100100110110010111000;
11'd920: out <= 32'b00001110110100110001001011000010;
11'd921: out <= 32'b00001100100110010000101001101100;
11'd922: out <= 32'b11110110101011001000010100001110;
11'd923: out <= 32'b10001001011100111111100100001011;
11'd924: out <= 32'b10100100100000110001110100000101;
11'd925: out <= 32'b01101001101101010101111000001001;
11'd926: out <= 32'b11010111111111011000001011100100;
11'd927: out <= 32'b10100000010101010101011110011110;
11'd928: out <= 32'b00110100111111011110011111110101;
11'd929: out <= 32'b11101101011110100111111110001100;
11'd930: out <= 32'b11111000110010110100100011111110;
11'd931: out <= 32'b00010010001001001101100111110001;
11'd932: out <= 32'b10011100011101010101000111011011;
11'd933: out <= 32'b00000001000101001000110100010100;
11'd934: out <= 32'b01000000010001100101010011110101;
11'd935: out <= 32'b01000101110110100110001111001111;
11'd936: out <= 32'b00010110011101101010110101111011;
11'd937: out <= 32'b11111100011000001010011110010101;
11'd938: out <= 32'b10001110110010010000001010000110;
11'd939: out <= 32'b00010010100010101000111010001001;
11'd940: out <= 32'b00001100101010011000110001111101;
11'd941: out <= 32'b00101000000001010000111100100100;
11'd942: out <= 32'b00100000011011011011000011100001;
11'd943: out <= 32'b11011101001111101111010011100111;
11'd944: out <= 32'b10101110010000101111011000000010;
11'd945: out <= 32'b11111001111000100010011101101101;
11'd946: out <= 32'b00110101011010111101010011110000;
11'd947: out <= 32'b00111110101101000010101010010101;
11'd948: out <= 32'b10011110101101010100111111001101;
11'd949: out <= 32'b10011100101111010111110101101001;
11'd950: out <= 32'b10010000101100111010111010010010;
11'd951: out <= 32'b11011011111010111110011110011001;
11'd952: out <= 32'b10010100111000100101010011110100;
11'd953: out <= 32'b01010111101001010001111111100101;
11'd954: out <= 32'b11110100001111001100001101101101;
11'd955: out <= 32'b11010111110110010000001011110110;
11'd956: out <= 32'b01110100101111100111010100000100;
11'd957: out <= 32'b00110111101100010010010001000101;
11'd958: out <= 32'b01010100011100100110010111110000;
11'd959: out <= 32'b11100000001011111100110100011000;
11'd960: out <= 32'b01000001000001100101101010110111;
11'd961: out <= 32'b00011001100111111000010101110111;
11'd962: out <= 32'b10011001111011000011000100011110;
11'd963: out <= 32'b10110111000011110000101101011001;
11'd964: out <= 32'b11011010010101110000101000000000;
11'd965: out <= 32'b10001000011001001101001001110010;
11'd966: out <= 32'b10100011000110010101111010110001;
11'd967: out <= 32'b01010111111111111000011110010010;
11'd968: out <= 32'b11110010001010011001011101001110;
11'd969: out <= 32'b11010101010111000001001000101101;
11'd970: out <= 32'b10100111101000111101011010101111;
11'd971: out <= 32'b11000100010000011000010010011111;
11'd972: out <= 32'b10011100001101010100100101000101;
11'd973: out <= 32'b11101100111011011011011000100010;
11'd974: out <= 32'b10001100110110111011100001000010;
11'd975: out <= 32'b10100010010101100100110011010011;
11'd976: out <= 32'b11111010001111100000100000110000;
11'd977: out <= 32'b11100111010110000100110010001010;
11'd978: out <= 32'b11000111101110110010111001100101;
11'd979: out <= 32'b01111010110100100100011111111000;
11'd980: out <= 32'b11101001110011100100010110000000;
11'd981: out <= 32'b01011101000000101010101001100010;
11'd982: out <= 32'b11100101100001010111010101101001;
11'd983: out <= 32'b00000000011010000011111010011000;
11'd984: out <= 32'b10110011110000011110110000010100;
11'd985: out <= 32'b00100010110100111010001000101111;
11'd986: out <= 32'b01110011011000100001111001100010;
11'd987: out <= 32'b11001100011001101110110001000010;
11'd988: out <= 32'b10101011010110000011110110100010;
11'd989: out <= 32'b01010111000110001110000100110011;
11'd990: out <= 32'b00000111000010110111001000000110;
11'd991: out <= 32'b10110110101101001110000100111001;
11'd992: out <= 32'b10001011001001000000001010111110;
11'd993: out <= 32'b11001111000011001101101100111110;
11'd994: out <= 32'b10001011001010011100101101110000;
11'd995: out <= 32'b10101001110011010110000110100010;
11'd996: out <= 32'b11010001000110100110011100110001;
11'd997: out <= 32'b11100001101001010111010011011001;
11'd998: out <= 32'b11111110111110100011101011010001;
11'd999: out <= 32'b00110111111001011111101100001111;
11'd1000: out <= 32'b01111001100111100101010001110110;
11'd1001: out <= 32'b01111011111011101101110101001111;
11'd1002: out <= 32'b01100110111001100101101100111101;
11'd1003: out <= 32'b10111001110000101101110010101001;
11'd1004: out <= 32'b01011101000000000011100000011010;
11'd1005: out <= 32'b00011101011001001011110110101110;
11'd1006: out <= 32'b11101011001010111000101111010111;
11'd1007: out <= 32'b11011100101010001001010000101111;
11'd1008: out <= 32'b00010000110101000011101110001101;
11'd1009: out <= 32'b00101010100111011110001100001100;
11'd1010: out <= 32'b11100000100000001010110000111000;
11'd1011: out <= 32'b11011011101001111111110101001111;
11'd1012: out <= 32'b00010111011101100111101011000100;
11'd1013: out <= 32'b01101011111010010111001100011111;
11'd1014: out <= 32'b01110010000001000110011001011011;
11'd1015: out <= 32'b00110011110001011111010011001110;
11'd1016: out <= 32'b11111100110010010011001111000100;
11'd1017: out <= 32'b10001111011100110101101110101000;
11'd1018: out <= 32'b11010011001001011101110010010011;
11'd1019: out <= 32'b00001011110100011110011011000111;
11'd1020: out <= 32'b00100001111101100110011101010011;
11'd1021: out <= 32'b01001110110011110110110000011110;
11'd1022: out <= 32'b10000011011011000001010001111010;
11'd1023: out <= 32'b11000000101000111100100110111010;
11'd1024: out <= 32'b10111001000011100111011010110111;
11'd1025: out <= 32'b00011101100001100011010111111100;
11'd1026: out <= 32'b10011101001011010001110111111101;
11'd1027: out <= 32'b01110101110111100100101001001101;
11'd1028: out <= 32'b10110010110101111011011010100010;
11'd1029: out <= 32'b10010001110001101111010001111010;
11'd1030: out <= 32'b00010001100101101010001101101111;
11'd1031: out <= 32'b10010100010011100100100011001001;
11'd1032: out <= 32'b01101110010110011111010110000010;
11'd1033: out <= 32'b01010010000111001101011111010000;
11'd1034: out <= 32'b10101010001011110011101010011010;
11'd1035: out <= 32'b01111110100000101101110100100110;
11'd1036: out <= 32'b10001001111001010011111001110010;
11'd1037: out <= 32'b11010011111011001010111111001101;
11'd1038: out <= 32'b11000010111100011000010100001100;
11'd1039: out <= 32'b01010011010011000011010100010001;
11'd1040: out <= 32'b01011001010011000101111010010110;
11'd1041: out <= 32'b10011110111100111111111111101010;
11'd1042: out <= 32'b01000011001110100110000100100101;
11'd1043: out <= 32'b00011010100010000110000011000011;
11'd1044: out <= 32'b10110111101101101101100001111100;
11'd1045: out <= 32'b01100111000001111010001010001000;
11'd1046: out <= 32'b11011001000010110000110110111011;
11'd1047: out <= 32'b11101010011011111100110110110010;
11'd1048: out <= 32'b10000000000110100010101101110000;
11'd1049: out <= 32'b11011010000111101001111111101101;
11'd1050: out <= 32'b10101101000110010011110111100011;
11'd1051: out <= 32'b11000011000011111100000001110001;
11'd1052: out <= 32'b01111111010101010001100111100111;
11'd1053: out <= 32'b10100010100000000101011111111010;
11'd1054: out <= 32'b00001100101100000111100101111111;
11'd1055: out <= 32'b00000010101001000010001110001001;
11'd1056: out <= 32'b00001101100100111011111010100010;
11'd1057: out <= 32'b01000001001010000111110010010011;
11'd1058: out <= 32'b11101011111011110010111011000101;
11'd1059: out <= 32'b10000110101110010001010110010000;
11'd1060: out <= 32'b01000001011010010101010110101011;
11'd1061: out <= 32'b01010110100011110101001100011000;
11'd1062: out <= 32'b11101111010000101010110110011011;
11'd1063: out <= 32'b11001011111100100001101011110010;
11'd1064: out <= 32'b01010101010100111110011110100000;
11'd1065: out <= 32'b10011001100101000011100111110100;
11'd1066: out <= 32'b00101111001010111000011111011010;
11'd1067: out <= 32'b01011000100010100101011001011101;
11'd1068: out <= 32'b00000010010010010001010010011010;
11'd1069: out <= 32'b11011100100001010100001000010110;
11'd1070: out <= 32'b10101100101100010001100000010111;
11'd1071: out <= 32'b00100111100011101010001011000100;
11'd1072: out <= 32'b00100100100011000101010010100110;
11'd1073: out <= 32'b11100010100010101110011111100001;
11'd1074: out <= 32'b10011111110101100101011111110000;
11'd1075: out <= 32'b00100111010000010010100111010100;
11'd1076: out <= 32'b11111000110010000110001000111101;
11'd1077: out <= 32'b11100101110100010000110100000100;
11'd1078: out <= 32'b10010010101011110010111111110101;
11'd1079: out <= 32'b00100001010111001111111111111001;
11'd1080: out <= 32'b01110100011011011100000001101110;
11'd1081: out <= 32'b00100101001101001010011001101011;
11'd1082: out <= 32'b01011110100000011111011011001000;
11'd1083: out <= 32'b11100111001100010011010001111111;
11'd1084: out <= 32'b10100100100110001011110100101000;
11'd1085: out <= 32'b00101101001000101000000100010010;
11'd1086: out <= 32'b00001000101000110111101000101111;
11'd1087: out <= 32'b00010111110100101001110010111100;
11'd1088: out <= 32'b10101000011101000001010111000001;
11'd1089: out <= 32'b11110110000110110100011110110011;
11'd1090: out <= 32'b10000101101000010110101000111001;
11'd1091: out <= 32'b11100001000101111111011111011010;
11'd1092: out <= 32'b11101110000111011000111001010110;
11'd1093: out <= 32'b00100100101111011010110111100011;
11'd1094: out <= 32'b11011111101100110000101010011110;
11'd1095: out <= 32'b10110101010011001100101101010101;
11'd1096: out <= 32'b11110011110001010101000001100001;
11'd1097: out <= 32'b01100001011011000101010100110010;
11'd1098: out <= 32'b11000010001001101111000011100010;
11'd1099: out <= 32'b00101000110000110101000001101110;
11'd1100: out <= 32'b11101001111001010100110101011100;
11'd1101: out <= 32'b11010110110110100110011110110101;
11'd1102: out <= 32'b00010011110101111101001100010111;
11'd1103: out <= 32'b11010100111000111110110111100111;
11'd1104: out <= 32'b10101110001001010111110111011101;
11'd1105: out <= 32'b11111111111011000101101101101000;
11'd1106: out <= 32'b11011000110110101001011000011010;
11'd1107: out <= 32'b01000111000110010110000001001010;
11'd1108: out <= 32'b11010110011001001001001001111111;
11'd1109: out <= 32'b10010001000100010000100101100001;
11'd1110: out <= 32'b10101001101000101000001010011001;
11'd1111: out <= 32'b10010101011100000000101000000010;
11'd1112: out <= 32'b01011111101100101100100000101100;
11'd1113: out <= 32'b01101100101010100101011110010011;
11'd1114: out <= 32'b01010001010010100111001000111011;
11'd1115: out <= 32'b10010010001111011111010011101010;
11'd1116: out <= 32'b00001101111001010110011100100111;
11'd1117: out <= 32'b01000101001110100001101101101010;
11'd1118: out <= 32'b01010101010001110001011001110101;
11'd1119: out <= 32'b10010100110110011011000001000010;
11'd1120: out <= 32'b11100100111101111000011111111111;
11'd1121: out <= 32'b00111011101101011001101010011011;
11'd1122: out <= 32'b10000100100110101010111101111111;
11'd1123: out <= 32'b00000111100010001111001010101100;
11'd1124: out <= 32'b10101100111110010001110000100111;
11'd1125: out <= 32'b10001010101110111110110011111000;
11'd1126: out <= 32'b11011010001100011000010001100010;
11'd1127: out <= 32'b01011000110001011000011011011001;
11'd1128: out <= 32'b01000000011101110001100100101111;
11'd1129: out <= 32'b10100010111110010011111110011011;
11'd1130: out <= 32'b01010011010110000011001001111001;
11'd1131: out <= 32'b10001110100100010011001000000011;
11'd1132: out <= 32'b00010111110100100010101111011100;
11'd1133: out <= 32'b10001000000010001100101101010100;
11'd1134: out <= 32'b10101001001100000100000101000101;
11'd1135: out <= 32'b00101000001001010110100010000111;
11'd1136: out <= 32'b00001101011001111100001100000101;
11'd1137: out <= 32'b01010001110011101110000000101110;
11'd1138: out <= 32'b01001111011000100010010010010001;
11'd1139: out <= 32'b01000010011010001011001111111000;
11'd1140: out <= 32'b00100111110011100011100111010010;
11'd1141: out <= 32'b11000011001001101111110110100101;
11'd1142: out <= 32'b01001111001100111000111000000010;
11'd1143: out <= 32'b01100110111101100000011011101011;
11'd1144: out <= 32'b00100011011000011101101101001011;
11'd1145: out <= 32'b10010010111011011011101000001011;
11'd1146: out <= 32'b00011011110000111111110101110101;
11'd1147: out <= 32'b11001100111001101110000100010010;
11'd1148: out <= 32'b00000110100001011011111001001010;
11'd1149: out <= 32'b01100101011111010010000000100011;
11'd1150: out <= 32'b10100000110011111101100011000101;
11'd1151: out <= 32'b10110010011111011010011110111111;
11'd1152: out <= 32'b01011110010110000101011110111100;
11'd1153: out <= 32'b01100110000100111100101110011001;
11'd1154: out <= 32'b11111111111100101010111111101011;
11'd1155: out <= 32'b00111100001010001101001001111110;
11'd1156: out <= 32'b00011110101001001010100001111001;
11'd1157: out <= 32'b10101010000001010111001111000101;
11'd1158: out <= 32'b00010011011010001111000000011011;
11'd1159: out <= 32'b00100100001000010011010110001010;
11'd1160: out <= 32'b11001000110001011010110111110110;
11'd1161: out <= 32'b11001001100111100111110001010000;
11'd1162: out <= 32'b01000111111110000111001000100011;
11'd1163: out <= 32'b00010011000101000001011110110110;
11'd1164: out <= 32'b10101111011100101100000100001010;
11'd1165: out <= 32'b11110101011101111001111110010100;
11'd1166: out <= 32'b10010000010101100110101000111010;
11'd1167: out <= 32'b00101010011000101010000100101110;
11'd1168: out <= 32'b00000000100110000010111111001101;
11'd1169: out <= 32'b01110000001011100010000001100000;
11'd1170: out <= 32'b11110111011011011011011000001100;
11'd1171: out <= 32'b10100010010110001011111111010011;
11'd1172: out <= 32'b10111101010010000001111000010011;
11'd1173: out <= 32'b00011000010110100111110101000001;
11'd1174: out <= 32'b10010110010010100101000000110100;
11'd1175: out <= 32'b11001100000001001000110010001101;
11'd1176: out <= 32'b11001000101100011101101101101100;
11'd1177: out <= 32'b00110101101010000100000110000010;
11'd1178: out <= 32'b10110011010010011111101110100000;
11'd1179: out <= 32'b01000001011010000011111110110111;
11'd1180: out <= 32'b11111100011101101000001110000110;
11'd1181: out <= 32'b11100100111000010100100101010100;
11'd1182: out <= 32'b00100001011101110011001110111101;
11'd1183: out <= 32'b10110100011100110011110111001011;
11'd1184: out <= 32'b01110100000110000010010101101110;
11'd1185: out <= 32'b11010100100010000011011100010001;
11'd1186: out <= 32'b11110010001111010000011011001001;
11'd1187: out <= 32'b01001001100011000010110111110011;
11'd1188: out <= 32'b00100111001010110000111010011010;
11'd1189: out <= 32'b11100010011001101000010110110011;
11'd1190: out <= 32'b00010100000101110011110100101110;
11'd1191: out <= 32'b11010111011000011100000000010100;
11'd1192: out <= 32'b11110101010110100101111110101010;
11'd1193: out <= 32'b00110111110000000100011011110110;
11'd1194: out <= 32'b01000111111000001110011000110001;
11'd1195: out <= 32'b10010001100010000000010101010101;
11'd1196: out <= 32'b10000111111101001110101011000101;
11'd1197: out <= 32'b01101101000011110000101011100110;
11'd1198: out <= 32'b01011011101001111101010101001110;
11'd1199: out <= 32'b01011001110000100000101011001011;
11'd1200: out <= 32'b10111011111111000010000101111011;
11'd1201: out <= 32'b00001000001011101011111111001010;
11'd1202: out <= 32'b10110110100100001011001010111111;
11'd1203: out <= 32'b01010101011011110101010111111011;
11'd1204: out <= 32'b01001100111000111011001000111110;
11'd1205: out <= 32'b01010010111000111010010010001001;
11'd1206: out <= 32'b00011000010110110100100010111010;
11'd1207: out <= 32'b11000011011000011001100111010111;
11'd1208: out <= 32'b10100000100011111010100110111011;
11'd1209: out <= 32'b01000010010110101011100001111001;
11'd1210: out <= 32'b01000000010000111100110010111101;
11'd1211: out <= 32'b00001000011001110000100011010111;
11'd1212: out <= 32'b01100100101101110011111111100111;
11'd1213: out <= 32'b00101001111111010010111110110001;
11'd1214: out <= 32'b00111111110011010110001111111111;
11'd1215: out <= 32'b00100001000000001010111111011011;
11'd1216: out <= 32'b10101010000110101101010000110000;
11'd1217: out <= 32'b01111110101111100111010011101111;
11'd1218: out <= 32'b01001111111000011010001011110010;
11'd1219: out <= 32'b11111011010000100010010011100011;
11'd1220: out <= 32'b10100110011111111011000001001011;
11'd1221: out <= 32'b00110111111100010010001100010011;
11'd1222: out <= 32'b10000001011011101000000100110011;
11'd1223: out <= 32'b10000100011010111110101100000100;
11'd1224: out <= 32'b01010101111010011000010101100110;
11'd1225: out <= 32'b00100010110110011011100011101111;
11'd1226: out <= 32'b00111101100010001111010000101100;
11'd1227: out <= 32'b11011100000100110000100001110000;
11'd1228: out <= 32'b00011010010000011000001110101110;
11'd1229: out <= 32'b01010101001000110010111010011010;
11'd1230: out <= 32'b01010010100000110101001100110110;
11'd1231: out <= 32'b11100111111001011111001011000011;
11'd1232: out <= 32'b11111011101100010101111011101010;
11'd1233: out <= 32'b01111011001101001010011000011011;
11'd1234: out <= 32'b11100000011011110011111111100111;
11'd1235: out <= 32'b01000101110011101000000100001110;
11'd1236: out <= 32'b01001100011101011001101010000000;
11'd1237: out <= 32'b11110001101011110011100001011101;
11'd1238: out <= 32'b01010110010000001010011010100011;
11'd1239: out <= 32'b01101010110010011010101111001110;
11'd1240: out <= 32'b01111111010001100111110111111110;
11'd1241: out <= 32'b01010001111011011111101111001010;
11'd1242: out <= 32'b00101010011011011011011100001100;
11'd1243: out <= 32'b10010100010110011100101100000100;
11'd1244: out <= 32'b00000100101011110001011001010110;
11'd1245: out <= 32'b01110101010101100001000111001101;
11'd1246: out <= 32'b11110010010011000001110101110000;
11'd1247: out <= 32'b10110111110111101000010101111100;
11'd1248: out <= 32'b00100010111101100100111011011011;
11'd1249: out <= 32'b10111000010001111110010010001101;
11'd1250: out <= 32'b11101000110010111001100101110100;
11'd1251: out <= 32'b01010111100011110100110111101011;
11'd1252: out <= 32'b10011011101000101111011101110101;
11'd1253: out <= 32'b11011111011010111100011011011100;
11'd1254: out <= 32'b11011010111010001011110011100100;
11'd1255: out <= 32'b11100011011111100000001011011001;
11'd1256: out <= 32'b10011100011011010000111010100000;
11'd1257: out <= 32'b10101110110001001011101010011110;
11'd1258: out <= 32'b10100100100001100000001110000100;
11'd1259: out <= 32'b01011100001001111011000011011110;
11'd1260: out <= 32'b11100001011101110100101001001100;
11'd1261: out <= 32'b11000000011110010111100110100010;
11'd1262: out <= 32'b01101001011000000001011101100000;
11'd1263: out <= 32'b10001011110000000011100100011100;
11'd1264: out <= 32'b11101001111100011110110100111010;
11'd1265: out <= 32'b11010111100001000101110010011010;
11'd1266: out <= 32'b00101111111001001000100000011110;
11'd1267: out <= 32'b10111101000010110100101100110010;
11'd1268: out <= 32'b11101101101001100000010011100000;
11'd1269: out <= 32'b11010101001101010011111110011010;
11'd1270: out <= 32'b11001101001101010011110001010010;
11'd1271: out <= 32'b01011011110000110010110000111010;
11'd1272: out <= 32'b11000111111000011010110001101101;
11'd1273: out <= 32'b00011111001110000111011010010011;
11'd1274: out <= 32'b10000001010001111100011010100100;
11'd1275: out <= 32'b01000110111001001110011000100100;
11'd1276: out <= 32'b01000100110100011001010000001110;
11'd1277: out <= 32'b01001000001010111100111001001011;
11'd1278: out <= 32'b01001111010100101101101101101000;
11'd1279: out <= 32'b10000100100001000110111001000100;
11'd1280: out <= 32'b11001011010001010001100000111000;
11'd1281: out <= 32'b10001101000111101001010010011110;
11'd1282: out <= 32'b10001010111110101010100111101010;
11'd1283: out <= 32'b10100000001111100111100101111001;
11'd1284: out <= 32'b11110011010001100100000100000011;
11'd1285: out <= 32'b11101000100111001001001010010010;
11'd1286: out <= 32'b11000000001001011001010011000111;
11'd1287: out <= 32'b11001000100000111110100100111011;
11'd1288: out <= 32'b10001101011001010101001011100011;
11'd1289: out <= 32'b11101100111110111110110101011001;
11'd1290: out <= 32'b00111100010101010100100110101011;
11'd1291: out <= 32'b10101101001110111011101101011011;
11'd1292: out <= 32'b00100000000000110101000010111001;
11'd1293: out <= 32'b01110100010001110011000111110100;
11'd1294: out <= 32'b11100110110101010100110111111111;
11'd1295: out <= 32'b01001011011010001100001010010101;
11'd1296: out <= 32'b01001101110010010011100011010000;
11'd1297: out <= 32'b10100001100010111101110010000111;
11'd1298: out <= 32'b01000110010101001100010000110101;
11'd1299: out <= 32'b01010110001110100000100010001100;
11'd1300: out <= 32'b11100011111010001111011011111011;
11'd1301: out <= 32'b11101101101000011100111100000110;
11'd1302: out <= 32'b00010011000111110010001111001010;
11'd1303: out <= 32'b01101111010000110101101100011101;
11'd1304: out <= 32'b01010011101001110101011010011111;
11'd1305: out <= 32'b01110000010100110101111000001110;
11'd1306: out <= 32'b10100001010011100100101111010101;
11'd1307: out <= 32'b10000110100100100000100000001101;
11'd1308: out <= 32'b11010100111010000110110111011010;
11'd1309: out <= 32'b00100011011100100011011100000001;
11'd1310: out <= 32'b01100101111101101011100001110110;
11'd1311: out <= 32'b00111011101110011010001010011101;
11'd1312: out <= 32'b11110000011100111000011111100010;
11'd1313: out <= 32'b01110000111111111000000111010101;
11'd1314: out <= 32'b10001011100111110001001001010000;
11'd1315: out <= 32'b10110100001010111001111110001001;
11'd1316: out <= 32'b10111010010010100110111100110000;
11'd1317: out <= 32'b01000010101000011001110011001101;
11'd1318: out <= 32'b10111010110001010011111111001000;
11'd1319: out <= 32'b11101110111011000000111110011001;
11'd1320: out <= 32'b01011100011010111100100101111101;
11'd1321: out <= 32'b10101000101111010110010000110000;
11'd1322: out <= 32'b10111111001000001010101011001010;
11'd1323: out <= 32'b11110001100000110101111011110001;
11'd1324: out <= 32'b00101110001010110010110010100001;
11'd1325: out <= 32'b01011000011110001001010111100001;
11'd1326: out <= 32'b10010111111110111000111100101111;
11'd1327: out <= 32'b11100110111101010110111111011110;
11'd1328: out <= 32'b01010011101000000000000010111111;
11'd1329: out <= 32'b01000111001101111101110011011110;
11'd1330: out <= 32'b11000100110111111000101010101010;
11'd1331: out <= 32'b11101110011001100110110000000011;
11'd1332: out <= 32'b11000000111101101110011110100100;
11'd1333: out <= 32'b11101110111010011010010000100111;
11'd1334: out <= 32'b11101001011011100001111011011100;
11'd1335: out <= 32'b01001101110000001001101000111100;
11'd1336: out <= 32'b11110010111100101000011011101100;
11'd1337: out <= 32'b00111001111101101001000000111110;
11'd1338: out <= 32'b11010111100010110101001101110110;
11'd1339: out <= 32'b11001000010111001000100011100100;
11'd1340: out <= 32'b00111010110010100001110110111100;
11'd1341: out <= 32'b01101110101010000111001101000001;
11'd1342: out <= 32'b00001000011110111110101001010011;
11'd1343: out <= 32'b01011101110010010101111001100001;
11'd1344: out <= 32'b10000110100001101100000000010101;
11'd1345: out <= 32'b00110001011111000000011110010111;
11'd1346: out <= 32'b01101010000011001000001010110101;
11'd1347: out <= 32'b11010000011000111010100111010101;
11'd1348: out <= 32'b00011011110001011010110110010000;
11'd1349: out <= 32'b11101011111100001011100111001001;
11'd1350: out <= 32'b00010101100001110111000111010010;
11'd1351: out <= 32'b01110101111101110010011001101101;
11'd1352: out <= 32'b00110111001010000001111001100111;
11'd1353: out <= 32'b00001110011010110100110001101110;
11'd1354: out <= 32'b00000111001001001110000100001111;
11'd1355: out <= 32'b10011001100101011000010101001010;
11'd1356: out <= 32'b10000001001010111111100111011111;
11'd1357: out <= 32'b11000000011101111011111100010001;
11'd1358: out <= 32'b01101111111011111100111001010001;
11'd1359: out <= 32'b10001100100101101000000010001000;
11'd1360: out <= 32'b11001101111010010111011110111111;
11'd1361: out <= 32'b10011110110110000100101101001011;
11'd1362: out <= 32'b11101111000110010111101100101110;
11'd1363: out <= 32'b10000110111011000011100001110011;
11'd1364: out <= 32'b01101011010001000001010111000010;
11'd1365: out <= 32'b01101111001100000110010010100010;
11'd1366: out <= 32'b00011011011000001110100011011100;
11'd1367: out <= 32'b00001011010011000001100100000100;
11'd1368: out <= 32'b10110100111111001110011110110001;
11'd1369: out <= 32'b01001010111101000101000010100010;
11'd1370: out <= 32'b00001111111000110110101010011111;
11'd1371: out <= 32'b01001011111010111110111111111010;
11'd1372: out <= 32'b00100010100111100110100010010111;
11'd1373: out <= 32'b10110000000001000001000110101100;
11'd1374: out <= 32'b01110111111010010010010110010100;
11'd1375: out <= 32'b00011011101101101010110011011101;
11'd1376: out <= 32'b00101100000001100111011010010000;
11'd1377: out <= 32'b01111010011100111110011010111011;
11'd1378: out <= 32'b01110111011101001000010011111000;
11'd1379: out <= 32'b10101000111011011001011101011010;
11'd1380: out <= 32'b10101111011100000010001111101101;
11'd1381: out <= 32'b11010010110011000011110000100011;
11'd1382: out <= 32'b11000100001111011100101010110011;
11'd1383: out <= 32'b00001110001101101011010000100101;
11'd1384: out <= 32'b00011011001110110111001010111001;
11'd1385: out <= 32'b00110100101010010011011010011000;
11'd1386: out <= 32'b11000000010100011001100110011011;
11'd1387: out <= 32'b00110011011101111000000100011101;
11'd1388: out <= 32'b00111111000010110001111010110111;
11'd1389: out <= 32'b01011101000001111001100101111100;
11'd1390: out <= 32'b00100010010110011010100110111010;
11'd1391: out <= 32'b10100110010011100110001100011111;
11'd1392: out <= 32'b00011011000111111111010001101000;
11'd1393: out <= 32'b01100100111000011000110101110001;
11'd1394: out <= 32'b01000011101000011110001110011101;
11'd1395: out <= 32'b10010110100010110111010111101010;
11'd1396: out <= 32'b10001111101000011000000110101100;
11'd1397: out <= 32'b01010000101001100111111010100100;
11'd1398: out <= 32'b11000110101101000010010000101111;
11'd1399: out <= 32'b00110111010000000001101001010000;
11'd1400: out <= 32'b00001000001101001001011011101010;
11'd1401: out <= 32'b11010100011011001100101111111000;
11'd1402: out <= 32'b01001011111001100111000001111001;
11'd1403: out <= 32'b11101110010011110101011101011111;
11'd1404: out <= 32'b01001111011111111110011000000110;
11'd1405: out <= 32'b01010010001011011100010010000011;
11'd1406: out <= 32'b10000100011011110010101010011110;
11'd1407: out <= 32'b00111000011110100011011111001001;
11'd1408: out <= 32'b10111010000101000110111001101110;
11'd1409: out <= 32'b01000100100100110010100111111110;
11'd1410: out <= 32'b00100001001001101111101111010100;
11'd1411: out <= 32'b00000010101010011001010010111100;
11'd1412: out <= 32'b01011100110010101100111010011011;
11'd1413: out <= 32'b00000001101001000100110101001101;
11'd1414: out <= 32'b01110110001111001010001100011001;
11'd1415: out <= 32'b10111100010001111010010110100000;
11'd1416: out <= 32'b00101111000101000010010111110001;
11'd1417: out <= 32'b00100101000110000111111100111001;
11'd1418: out <= 32'b10010001100000011110011001100111;
11'd1419: out <= 32'b01101111001100111000110101001011;
11'd1420: out <= 32'b10100111010101011101110101101011;
11'd1421: out <= 32'b11111101001100100000110111011001;
11'd1422: out <= 32'b10100100111101001010111100000000;
11'd1423: out <= 32'b11001000011110101111010000011100;
11'd1424: out <= 32'b11101011101100110100111100010111;
11'd1425: out <= 32'b10110011011100101010011100110000;
11'd1426: out <= 32'b00110100001010000010011011010010;
11'd1427: out <= 32'b00001110011111111010010011000110;
11'd1428: out <= 32'b11110111111010101111001110100011;
11'd1429: out <= 32'b11100101100010110101101100111010;
11'd1430: out <= 32'b10001100001111011100001011110101;
11'd1431: out <= 32'b01100110101000110000111011000101;
11'd1432: out <= 32'b01101010010101111001001111000101;
11'd1433: out <= 32'b01111001010011011110101111001100;
11'd1434: out <= 32'b10101000000011010111101101100110;
11'd1435: out <= 32'b10011011110011000110000110000001;
11'd1436: out <= 32'b11001000101100100011000110100000;
11'd1437: out <= 32'b01011101110001101001000110011001;
11'd1438: out <= 32'b11100100100010001010001001110010;
11'd1439: out <= 32'b00010011100111101010110101110001;
11'd1440: out <= 32'b01110100100010010000011100111110;
11'd1441: out <= 32'b01000110010011010011110010111110;
11'd1442: out <= 32'b10011100000110111010100111001101;
11'd1443: out <= 32'b01010000101110111011110111101011;
11'd1444: out <= 32'b00101111100101000011110110101001;
11'd1445: out <= 32'b00110011101100001110110011100000;
11'd1446: out <= 32'b10100011010010001000110111111011;
11'd1447: out <= 32'b01110101101111000000011101010001;
11'd1448: out <= 32'b01100100011001110110111101001011;
11'd1449: out <= 32'b00100001000001010100001001111011;
11'd1450: out <= 32'b10100010110111010101110100011111;
11'd1451: out <= 32'b00111100110110000110001010110000;
11'd1452: out <= 32'b01111011001101001110001001110001;
11'd1453: out <= 32'b00011011100001101100010101010110;
11'd1454: out <= 32'b00101001011001011010001010010000;
11'd1455: out <= 32'b11101101000111111100010000010001;
11'd1456: out <= 32'b11000110000111111011001001100000;
11'd1457: out <= 32'b10101000011111011001111110110001;
11'd1458: out <= 32'b00011001000001011100111011000111;
11'd1459: out <= 32'b11100100010010101110101010110011;
11'd1460: out <= 32'b11001000110010001000111011001000;
11'd1461: out <= 32'b11000110000101110000111011101100;
11'd1462: out <= 32'b01000101000100101010110111111000;
11'd1463: out <= 32'b00000100010100000111110000100011;
11'd1464: out <= 32'b10010010011000110000011101001010;
11'd1465: out <= 32'b01011110011100010010111001011010;
11'd1466: out <= 32'b10011001111010010011101110110101;
11'd1467: out <= 32'b10001011001011011011110011111000;
11'd1468: out <= 32'b11011100010111111110001001100111;
11'd1469: out <= 32'b01111110110110001000010010011011;
11'd1470: out <= 32'b11001010100001110010111111110011;
11'd1471: out <= 32'b10011001011010111111101011101010;
11'd1472: out <= 32'b10011100000000011111010000011110;
11'd1473: out <= 32'b10011011010001001011011100111001;
11'd1474: out <= 32'b11101011010010110000110001111110;
11'd1475: out <= 32'b10001000000001000001010010110101;
11'd1476: out <= 32'b01100111100010010011010110111110;
11'd1477: out <= 32'b10000110011101000010000101010100;
11'd1478: out <= 32'b01010101111110110000010111000111;
11'd1479: out <= 32'b10110010010010001111001101001011;
11'd1480: out <= 32'b01010110001001101100101101110100;
11'd1481: out <= 32'b10100101101000101011110101101000;
11'd1482: out <= 32'b01110010001001100010001101010000;
11'd1483: out <= 32'b01010100010001000110001010000011;
11'd1484: out <= 32'b00000111110110111110100010110110;
11'd1485: out <= 32'b01110001110100110011000101011101;
11'd1486: out <= 32'b01001101001100100010110000011111;
11'd1487: out <= 32'b11011111100100110010001110011110;
11'd1488: out <= 32'b01011111011111111111011010001010;
11'd1489: out <= 32'b10101100110100011100110011111000;
11'd1490: out <= 32'b01001111010110110111010111010000;
11'd1491: out <= 32'b10010011000000110110011101100010;
11'd1492: out <= 32'b10011101001110101110111011001010;
11'd1493: out <= 32'b01011001101010100100110100110100;
11'd1494: out <= 32'b00101111010101011001010010010010;
11'd1495: out <= 32'b10010000011110110000101001101100;
11'd1496: out <= 32'b00010011000000111000001001010101;
11'd1497: out <= 32'b11110001011000111010100001100011;
11'd1498: out <= 32'b11100111100011101010001101000111;
11'd1499: out <= 32'b10011010000110000100011110010110;
11'd1500: out <= 32'b00010111001001110101111111100000;
11'd1501: out <= 32'b00000100000110100100101110000010;
11'd1502: out <= 32'b01000111111101111100111101101111;
11'd1503: out <= 32'b01100011000000100010000000101101;
11'd1504: out <= 32'b11111011011101010011101101111010;
11'd1505: out <= 32'b01011101111100000001101011111110;
11'd1506: out <= 32'b00001101001100010000111011100010;
11'd1507: out <= 32'b01110000001111011001110000101111;
11'd1508: out <= 32'b01111100100101011011010010001001;
11'd1509: out <= 32'b00011110010010110001100111000101;
11'd1510: out <= 32'b10010011011111011101011011101111;
11'd1511: out <= 32'b00001111110110111000111010101110;
11'd1512: out <= 32'b00100001100001000001111100110010;
11'd1513: out <= 32'b11110110101000011110001101101010;
11'd1514: out <= 32'b01010010000010000010010011001110;
11'd1515: out <= 32'b01111100001101100110110010000001;
11'd1516: out <= 32'b00111110111100110101000110001010;
11'd1517: out <= 32'b01011100010100101010110001000101;
11'd1518: out <= 32'b00001100000001011000111010000100;
11'd1519: out <= 32'b00001110100000111110000101100010;
11'd1520: out <= 32'b00111110111011000011101001010101;
11'd1521: out <= 32'b01011101100110101010001001100100;
11'd1522: out <= 32'b01010101001010110001001110100111;
11'd1523: out <= 32'b00110110100111001011001001111000;
11'd1524: out <= 32'b10101100111100101001111111100101;
11'd1525: out <= 32'b01110100100001010101110101010101;
11'd1526: out <= 32'b00111000100100100010111101001001;
11'd1527: out <= 32'b01010011110101000000001011011000;
11'd1528: out <= 32'b00111011111101000000101001100011;
11'd1529: out <= 32'b00110000110000010010111101101101;
11'd1530: out <= 32'b00001010101101111001000001010010;
11'd1531: out <= 32'b10100110010001110000011101001100;
11'd1532: out <= 32'b11001010110101111110101101110001;
11'd1533: out <= 32'b10110010100101101000110011000010;
11'd1534: out <= 32'b11011111111001101111111001100110;
11'd1535: out <= 32'b10100000001111110010000001011100;
11'd1536: out <= 32'b01111001110100101010101100110100;
11'd1537: out <= 32'b10010000100110010000010110001110;
11'd1538: out <= 32'b01010010011000111011111110011100;
11'd1539: out <= 32'b10111001111011001111100100110010;
11'd1540: out <= 32'b11111101010100011010100111000011;
11'd1541: out <= 32'b00100100110101000001010011011001;
11'd1542: out <= 32'b11110011101001111100010110101010;
11'd1543: out <= 32'b00110011110111010101011001111011;
11'd1544: out <= 32'b11010001011110101000101010000001;
11'd1545: out <= 32'b00110111101000010111000101100111;
11'd1546: out <= 32'b10001101111101011010111111110101;
11'd1547: out <= 32'b00001100101001001011001010100100;
11'd1548: out <= 32'b10101100111101101110000101001111;
11'd1549: out <= 32'b01100011100000011110010010001101;
11'd1550: out <= 32'b01101011010001001101110000001111;
11'd1551: out <= 32'b11011001111011101001101000011011;
11'd1552: out <= 32'b01101001010101111010111001001101;
11'd1553: out <= 32'b10111100101000110111000100101010;
11'd1554: out <= 32'b11001111010000011000011011010000;
11'd1555: out <= 32'b01010100011011010101001011010110;
11'd1556: out <= 32'b11111010010100100100111100100101;
11'd1557: out <= 32'b10010100011101000110011010011001;
11'd1558: out <= 32'b01110001011100111111001101100110;
11'd1559: out <= 32'b01111110110000111001001111010110;
11'd1560: out <= 32'b10010011101100110101001001101010;
11'd1561: out <= 32'b01101001101101101010100000011001;
11'd1562: out <= 32'b11000101001101111100111001110000;
11'd1563: out <= 32'b00011000100110100101000110100001;
11'd1564: out <= 32'b11111111000000100010101010000101;
11'd1565: out <= 32'b10100010000110001111001101101010;
11'd1566: out <= 32'b10001100100110011101000111101111;
11'd1567: out <= 32'b10000110100101001101000001000000;
11'd1568: out <= 32'b10001111001000000110000100100100;
11'd1569: out <= 32'b01101000111011101110001111101111;
11'd1570: out <= 32'b01011101011010000000001111010111;
11'd1571: out <= 32'b01111000101011010111101110101111;
11'd1572: out <= 32'b11111000010100110000000011111111;
11'd1573: out <= 32'b10110001111011100000100000011010;
11'd1574: out <= 32'b01001110101010010111000101101100;
11'd1575: out <= 32'b01101111110101111111100011001000;
11'd1576: out <= 32'b11101101010101001000011100111001;
11'd1577: out <= 32'b10010111100110110111110011010000;
11'd1578: out <= 32'b10010100110101111011100000010100;
11'd1579: out <= 32'b00111010110100000000101010001111;
11'd1580: out <= 32'b00111110100110110110010101111110;
11'd1581: out <= 32'b11000000001101100101010000101000;
11'd1582: out <= 32'b01110010010100000100001011101101;
11'd1583: out <= 32'b01000010101110100010100010010101;
11'd1584: out <= 32'b00010111010001011101101011010101;
11'd1585: out <= 32'b10111110100000010001000011110000;
11'd1586: out <= 32'b10100010000010110001101001010000;
11'd1587: out <= 32'b01010100000001011001111000000101;
11'd1588: out <= 32'b10000110110100101010101011110110;
11'd1589: out <= 32'b00110110001111110001001110110000;
11'd1590: out <= 32'b11100001001001011001011010001110;
11'd1591: out <= 32'b11101101111010001000010100111000;
11'd1592: out <= 32'b11000001101100100111111110101111;
11'd1593: out <= 32'b01001100110110001001001110111101;
11'd1594: out <= 32'b11001110001001000001111111111101;
11'd1595: out <= 32'b00001001011111000101111100111001;
11'd1596: out <= 32'b10111100001000000001010000100001;
11'd1597: out <= 32'b01000111010111010011101001010001;
11'd1598: out <= 32'b01000100101110100001010101100110;
11'd1599: out <= 32'b11010000111001011011001010011000;
11'd1600: out <= 32'b10101000101000011101010001011010;
11'd1601: out <= 32'b00011111101001100101010100100001;
11'd1602: out <= 32'b11101110100110001100000010000101;
11'd1603: out <= 32'b01111101000101110111101011110010;
11'd1604: out <= 32'b01101101011011011101001100001011;
11'd1605: out <= 32'b10010011101001011000110101100111;
11'd1606: out <= 32'b01011101010000100010010111000110;
11'd1607: out <= 32'b11110101101011111010101011011000;
11'd1608: out <= 32'b11101010010011001101100111011011;
11'd1609: out <= 32'b00101111000000110011111101011000;
11'd1610: out <= 32'b11010001000001000100100000011000;
11'd1611: out <= 32'b01011010100000001100111010000011;
11'd1612: out <= 32'b10010011010011001001010001011001;
11'd1613: out <= 32'b11000011100111001001100001010010;
11'd1614: out <= 32'b11110101111001001111111011001101;
11'd1615: out <= 32'b11000110011100011111101001011110;
11'd1616: out <= 32'b01000111101000111110011111001010;
11'd1617: out <= 32'b10011000110101111100011000111000;
11'd1618: out <= 32'b10000001010101010100100101011011;
11'd1619: out <= 32'b10111100111000000110000000010011;
11'd1620: out <= 32'b01000011000111100010000101100110;
11'd1621: out <= 32'b01000001111001100100000100011000;
11'd1622: out <= 32'b11010000110101010101010101000011;
11'd1623: out <= 32'b01000010001110001101000110110101;
11'd1624: out <= 32'b10110011010001001010100100011111;
11'd1625: out <= 32'b01111011111000011011001000110111;
11'd1626: out <= 32'b10001000110110001000011011111000;
11'd1627: out <= 32'b01110011011000010111000111111010;
11'd1628: out <= 32'b11111100011101100000101001101000;
11'd1629: out <= 32'b01111101100000011001100101000010;
11'd1630: out <= 32'b11110110100100001011111101100100;
11'd1631: out <= 32'b00001111001000010001110101110000;
11'd1632: out <= 32'b01111010010101000000010101010010;
11'd1633: out <= 32'b10100100110100110010001010011011;
11'd1634: out <= 32'b01000001100010100101110110101011;
11'd1635: out <= 32'b00110011000111110100000001100100;
11'd1636: out <= 32'b11000010111100101011111111110001;
11'd1637: out <= 32'b00110010111100001110010000010001;
11'd1638: out <= 32'b11001100001101000010110100111111;
11'd1639: out <= 32'b01000011011000101001000101010100;
11'd1640: out <= 32'b11001001110000100001100110011100;
11'd1641: out <= 32'b00001101111010110010111011111010;
11'd1642: out <= 32'b10001101111010111101111101100000;
11'd1643: out <= 32'b11101110001000000101100110111010;
11'd1644: out <= 32'b11001101000000010001110111111101;
11'd1645: out <= 32'b00111011011111100100000011000111;
11'd1646: out <= 32'b00001010000011000001100011111111;
11'd1647: out <= 32'b11001000111010100011100101001000;
11'd1648: out <= 32'b00010010100111111001010000011001;
11'd1649: out <= 32'b10110010000111011010011100110001;
11'd1650: out <= 32'b00001011010101100011111001101011;
11'd1651: out <= 32'b00001011110110100000100110101011;
11'd1652: out <= 32'b10110100111101001011001011100110;
11'd1653: out <= 32'b10010111100011100110101000100010;
11'd1654: out <= 32'b01100000110010011110010110110011;
11'd1655: out <= 32'b00001010001100011101101011010011;
11'd1656: out <= 32'b11101000011000111000000010011100;
11'd1657: out <= 32'b01111110111111001001111111000100;
11'd1658: out <= 32'b00110011100111100111101100001111;
11'd1659: out <= 32'b10101111010111011111101001000100;
11'd1660: out <= 32'b10111100111011111100100111101001;
11'd1661: out <= 32'b01011000001001000010010010110100;
11'd1662: out <= 32'b00111010111111000100001110010000;
11'd1663: out <= 32'b00001011101010010001111100011010;
11'd1664: out <= 32'b00000000000000010000000000111110;
11'd1665: out <= 32'b00000000000000110000000000000010;
11'd1666: out <= 32'b00000000000001010000000000000100;
11'd1667: out <= 32'b00000000000001110000000000000110;
11'd1668: out <= 32'b00000000000010010000000000001000;
11'd1669: out <= 32'b00000000000000010000000000001010;
11'd1670: out <= 32'b00000000000011110000000000000000;
11'd1671: out <= 32'b01101111000000101110011001010000;
11'd1672: out <= 32'b10010001101011001010101010010010;
11'd1673: out <= 32'b01000010101001010011111101101111;
11'd1674: out <= 32'b10011101100101110001110101101011;
11'd1675: out <= 32'b10110110110011001101100010000101;
11'd1676: out <= 32'b01011001110101011000001100101011;
11'd1677: out <= 32'b01100101111010011010010001110000;
11'd1678: out <= 32'b01111010010110000000101000110010;
11'd1679: out <= 32'b10001110110111101010011101101110;
11'd1680: out <= 32'b10011111110000111100000100111000;
11'd1681: out <= 32'b10100011110011000111010000011100;
11'd1682: out <= 32'b00001010011100001000000010101001;
11'd1683: out <= 32'b00110100110110100100100011010000;
11'd1684: out <= 32'b00110101111001110100010111010101;
11'd1685: out <= 32'b01111011000100000011001110000000;
11'd1686: out <= 32'b01101000101011010110100011110011;
11'd1687: out <= 32'b10001010000001001100000010101110;
11'd1688: out <= 32'b00010111101010001101010001100100;
11'd1689: out <= 32'b00110010101101101110001110110001;
11'd1690: out <= 32'b11100101100001011111011010101000;
11'd1691: out <= 32'b11111111110110010101111110110011;
11'd1692: out <= 32'b00111111100111100101011011101011;
11'd1693: out <= 32'b10101110110100111010001101111101;
11'd1694: out <= 32'b01000101010110110000100000110000;
11'd1695: out <= 32'b11111010110110110000011010111001;
11'd1696: out <= 32'b10100000011010010110011001110001;
11'd1697: out <= 32'b11011110011110100011110100100011;
11'd1698: out <= 32'b10000010010111010011100110010001;
11'd1699: out <= 32'b00101100010101000111011000001011;
11'd1700: out <= 32'b00110010100101010011100010001101;
11'd1701: out <= 32'b11110000111101110100100110011010;
11'd1702: out <= 32'b00111101101010111110011100111011;
11'd1703: out <= 32'b11100010011001000000010011011110;
11'd1704: out <= 32'b01111001000001111000001101001000;
11'd1705: out <= 32'b10010100111110111001111100110010;
11'd1706: out <= 32'b01010101110110111100000011010011;
11'd1707: out <= 32'b00110011110110000111011010011101;
11'd1708: out <= 32'b11101100111101101000001100010010;
11'd1709: out <= 32'b00101000010001011100101000000010;
11'd1710: out <= 32'b10101110111110000001010000110101;
11'd1711: out <= 32'b01110010111101100110110001100110;
11'd1712: out <= 32'b00111111000100010011001000011100;
11'd1713: out <= 32'b01010010011101100011101011100001;
11'd1714: out <= 32'b01101010111100000011100000001001;
11'd1715: out <= 32'b11000111010110001111110110111010;
11'd1716: out <= 32'b00000011101001111010110010100011;
11'd1717: out <= 32'b01000000100101111110100010101101;
11'd1718: out <= 32'b10001010100011000011000010111000;
11'd1719: out <= 32'b11000111100011101110001000101000;
11'd1720: out <= 32'b00110101000000000011110110011111;
11'd1721: out <= 32'b10000011111011101011101101011000;
11'd1722: out <= 32'b01000001010001111110101010110111;
11'd1723: out <= 32'b11100101000100001000010110000010;
11'd1724: out <= 32'b10001010001100101011100100010000;
11'd1725: out <= 32'b00110000011010000101010010101100;
11'd1726: out <= 32'b00010101010111001010000101011100;
11'd1727: out <= 32'b11100101111101011101111111001011;
11'd1728: out <= 32'b00011010010000100110101100110001;
11'd1729: out <= 32'b10100110111101000100111010111110;
11'd1730: out <= 32'b00010100111010010000010100000110;
11'd1731: out <= 32'b01011011111110000110101000010101;
11'd1732: out <= 32'b00100101001100101001111111011100;
11'd1733: out <= 32'b00100010100010000010010010100011;
11'd1734: out <= 32'b11010000101101000101011001011000;
11'd1735: out <= 32'b10000011000000001001011011000100;
11'd1736: out <= 32'b01000000001010100100101010000100;
11'd1737: out <= 32'b01000001101010001000010011010101;
11'd1738: out <= 32'b10101010101001010011101011100000;
11'd1739: out <= 32'b11100010001100111000100011010001;
11'd1740: out <= 32'b10000100101001100100010000011110;
11'd1741: out <= 32'b01001100110000001001110110011101;
11'd1742: out <= 32'b00000001010011101011011111101101;
11'd1743: out <= 32'b01010010011110101001111011011100;
11'd1744: out <= 32'b10100011110111000010001010110011;
11'd1745: out <= 32'b00100100000111000011011010010011;
11'd1746: out <= 32'b00110010100000001001001110001111;
11'd1747: out <= 32'b10101010111101110110001101101010;
11'd1748: out <= 32'b00110011101100001001000001110001;
11'd1749: out <= 32'b11111111101000110000010101000111;
11'd1750: out <= 32'b01100101010111010000010110110010;
11'd1751: out <= 32'b11110010010111011000110110101100;
11'd1752: out <= 32'b00000111011111011111001101010011;
11'd1753: out <= 32'b11100100001101100101101010000111;
11'd1754: out <= 32'b11000011100100010011010001000110;
11'd1755: out <= 32'b01101000101010110111111111111000;
11'd1756: out <= 32'b00101010100010010111100010011010;
11'd1757: out <= 32'b01011110000000101010010110110101;
11'd1758: out <= 32'b01111001110011101011001101110010;
11'd1759: out <= 32'b00111010000101101100100001010111;
11'd1760: out <= 32'b00101001100110000011101100110001;
11'd1761: out <= 32'b00101111110000100000011011000110;
11'd1762: out <= 32'b00110100001110001010001001111000;
11'd1763: out <= 32'b10010101100011110010011100000111;
11'd1764: out <= 32'b11001111110011100011001010000100;
11'd1765: out <= 32'b11110100101111101101011001110111;
11'd1766: out <= 32'b10110100011110000000110000010000;
11'd1767: out <= 32'b00111110111110000101110010110000;
11'd1768: out <= 32'b10111101001101111100010111100111;
11'd1769: out <= 32'b10100111110111100100011100111010;
11'd1770: out <= 32'b00101011110100101000110010110111;
11'd1771: out <= 32'b10110010001011000100100001111011;
11'd1772: out <= 32'b10101001101110100011100000011110;
11'd1773: out <= 32'b01000000110111001000110101010010;
11'd1774: out <= 32'b10001001010001011010101010101101;
11'd1775: out <= 32'b11001110000000111100010010100011;
11'd1776: out <= 32'b00011011011011101001000110101010;
11'd1777: out <= 32'b00110100101010001100011100101000;
11'd1778: out <= 32'b00000100010111010011011000001110;
11'd1779: out <= 32'b11101110001001001011011001111101;
11'd1780: out <= 32'b00111001111001001000110110100010;
11'd1781: out <= 32'b01000010100100101011011101001000;
11'd1782: out <= 32'b11000100011101010100010000110010;
11'd1783: out <= 32'b11010000001101100111011010110100;
11'd1784: out <= 32'b10100100101001110101110001101001;
11'd1785: out <= 32'b10100011100000110011111111011011;
11'd1786: out <= 32'b10010001100111111110001100010100;
11'd1787: out <= 32'b11001000111110001000010110111101;
11'd1788: out <= 32'b00011001101001000001001011101000;
11'd1789: out <= 32'b11111100101010001111000010111011;
11'd1790: out <= 32'b11100101110110110000010000111010;
11'd1791: out <= 32'b11000010111101001100001011110100;
11'd1792: out <= 32'b00000000000000000000000000000000;
11'd1793: out <= 32'b00000000000000000000000000000000;
11'd1794: out <= 32'b00000000000000000000000000000000;
11'd1795: out <= 32'b00000000000000000000000000000000;
11'd1796: out <= 32'b00000011110000000000000000000000;
11'd1797: out <= 32'b00110000000011000000110000110000;
11'd1798: out <= 32'b00001100001100000011000000001100;
11'd1799: out <= 32'b00000000000000000000001111000000;
11'd1800: out <= 32'b00000000111100000000000000000000;
11'd1801: out <= 32'b00001100001100000000001100110000;
11'd1802: out <= 32'b00000000001100000000000000110000;
11'd1803: out <= 32'b00000000000000000000000000110000;
11'd1804: out <= 32'b00000011111100000000000000000000;
11'd1805: out <= 32'b00000000000011000000110000001100;
11'd1806: out <= 32'b00000000110000000000000000110000;
11'd1807: out <= 32'b00000000000000000000111111111100;
11'd1808: out <= 32'b00001111111100000000000000000000;
11'd1809: out <= 32'b00000000000011000000000000001100;
11'd1810: out <= 32'b00000000000011000000001111110000;
11'd1811: out <= 32'b00000000000000000000111111110000;
11'd1812: out <= 32'b00000011000000000000000000000000;
11'd1813: out <= 32'b00110000110000000000110000000000;
11'd1814: out <= 32'b00000000110000000011111111110000;
11'd1815: out <= 32'b00000000000000000000000011000000;
11'd1816: out <= 32'b00111111111111000000000000000000;
11'd1817: out <= 32'b00110000000000000011000000000000;
11'd1818: out <= 32'b00000000000011000000111111111100;
11'd1819: out <= 32'b00000000000000000000111111110000;
11'd1820: out <= 32'b00000011111111000000000000000000;
11'd1821: out <= 32'b00110000000000000000110000000000;
11'd1822: out <= 32'b00110000000011000011111111110000;
11'd1823: out <= 32'b00000000000000000000111111110000;
11'd1824: out <= 32'b00111111111111000000000000000000;
11'd1825: out <= 32'b00000000001100000000000000001100;
11'd1826: out <= 32'b00000000110000000000000000110000;
11'd1827: out <= 32'b00000000000000000000001100000000;
11'd1828: out <= 32'b00001111111100000000000000000000;
11'd1829: out <= 32'b00110000000011000011000000001100;
11'd1830: out <= 32'b00110000000011000000111111110000;
11'd1831: out <= 32'b00000000000000000000111111110000;
11'd1832: out <= 32'b00001111111100000000000000000000;
11'd1833: out <= 32'b00110000000011000011000000001100;
11'd1834: out <= 32'b00000000000011000000111111111100;
11'd1835: out <= 32'b00000000000000000000111111110000;
11'd1836: out <= 32'b00000000000000000000000000000000;
11'd1837: out <= 32'b00000000000000000000000000000000;
11'd1838: out <= 32'b00000000000000000000111111110000;
11'd1839: out <= 32'b00000000000000000000000000000000;
11'd1840: out <= 32'b10011011011011100001000110110100;
11'd1841: out <= 32'b00010010011101000110111000101111;
11'd1842: out <= 32'b00011110110010001100010011100111;
11'd1843: out <= 32'b01101110101111111100011111100110;
11'd1844: out <= 32'b00011100001110011001000101001010;
11'd1845: out <= 32'b00010101000010010010111001000111;
11'd1846: out <= 32'b00000001010110000000101101100000;
11'd1847: out <= 32'b01001011110000101111101101001010;
11'd1848: out <= 32'b10110110010100111100010000010000;
11'd1849: out <= 32'b11100101101100010100011101000000;
11'd1850: out <= 32'b01101101100010100101111001111110;
11'd1851: out <= 32'b11000101100000101011110011000010;
11'd1852: out <= 32'b11001111100100001000000010111110;
11'd1853: out <= 32'b10110010100100011010000100011110;
11'd1854: out <= 32'b10100111011000011011100100111010;
11'd1855: out <= 32'b00010010101001011100000101111110;
11'd1856: out <= 32'b00111011011000000000000110110101;
11'd1857: out <= 32'b11101010010011010100010110110001;
11'd1858: out <= 32'b11011001010001101100101101010111;
11'd1859: out <= 32'b11011010011000011011101100010011;
11'd1860: out <= 32'b11001101111011010100011111111011;
11'd1861: out <= 32'b01100000100110001101000111010010;
11'd1862: out <= 32'b11000001010101101011011010010101;
11'd1863: out <= 32'b00000100011111001001111101101111;
11'd1864: out <= 32'b11000101011010110011111111011010;
11'd1865: out <= 32'b10011011101011001000111100000110;
11'd1866: out <= 32'b01110100011111100111011110100011;
11'd1867: out <= 32'b00110100101010000110011000111101;
11'd1868: out <= 32'b00111011101100011100001100001010;
11'd1869: out <= 32'b00011110110111101110000010001110;
11'd1870: out <= 32'b11011100110100000110100011000100;
11'd1871: out <= 32'b01001101111100000100110010001000;
11'd1872: out <= 32'b01011111001100000010011011011011;
11'd1873: out <= 32'b00011100001001010001110101110111;
11'd1874: out <= 32'b11000011010001011010011001010010;
11'd1875: out <= 32'b11100011010010101010011011010111;
11'd1876: out <= 32'b10011111110110111011100100000000;
11'd1877: out <= 32'b11100100100011110001111100000111;
11'd1878: out <= 32'b11011001010001011001001000110011;
11'd1879: out <= 32'b10101110000001011101110110101000;
11'd1880: out <= 32'b01111101001110011000011101110011;
11'd1881: out <= 32'b11001100001111001001111111111000;
11'd1882: out <= 32'b11110101010010110011001101101000;
11'd1883: out <= 32'b00100100111000100001000000000111;
11'd1884: out <= 32'b01101010100110100011010110101001;
11'd1885: out <= 32'b01011010001101101100110011010100;
11'd1886: out <= 32'b00011111100010000111001101111101;
11'd1887: out <= 32'b11011111111001000011001111000000;
11'd1888: out <= 32'b00011001100000001110111010010100;
11'd1889: out <= 32'b00010100010011010010100110011011;
11'd1890: out <= 32'b10110101100100111111100111111001;
11'd1891: out <= 32'b11011000010100001011000111001001;
11'd1892: out <= 32'b01001011110111001010111101000010;
11'd1893: out <= 32'b10111011111001111010000001000100;
11'd1894: out <= 32'b00110001011101000011111001100110;
11'd1895: out <= 32'b11101100110100011100000101000100;
11'd1896: out <= 32'b10101001000001101110011101110001;
11'd1897: out <= 32'b00000011111011001001011001111100;
11'd1898: out <= 32'b00110111101010010001111111010010;
11'd1899: out <= 32'b00001001011101010101100100001101;
11'd1900: out <= 32'b11011101111101010001110000010110;
11'd1901: out <= 32'b10010001101001111011100001110101;
11'd1902: out <= 32'b00110100000100100110111001101110;
11'd1903: out <= 32'b00000100011100101111001011011010;
11'd1904: out <= 32'b01001100010010000001000000001111;
11'd1905: out <= 32'b11010110010011001000100011101000;
11'd1906: out <= 32'b00101001000101101101001011000100;
11'd1907: out <= 32'b10010001111111101001101001100001;
11'd1908: out <= 32'b10001100001000111011000100010000;
11'd1909: out <= 32'b10001111111011100110010011100000;
11'd1910: out <= 32'b00111010000110000011110000110111;
11'd1911: out <= 32'b11100100000111111110000110001011;
11'd1912: out <= 32'b00001111111100000000000110000000;
11'd1913: out <= 32'b00110000000000000011000110001100;
11'd1914: out <= 32'b00000000000011000000111111110000;
11'd1915: out <= 32'b00000011000000000000111111110000;
11'd1916: out <= 32'b01111010101101110010010000100110;
11'd1917: out <= 32'b01110100011110011101010100010101;
11'd1918: out <= 32'b11011111111111100010101001100011;
11'd1919: out <= 32'b11001010011100100101000110000010;
11'd1920: out <= 32'b00001111000000000000000000000000;
11'd1921: out <= 32'b00110000000011000011000011110000;
11'd1922: out <= 32'b00110000000011000011111111111100;
11'd1923: out <= 32'b00000000000000000011000000001100;
11'd1924: out <= 32'b00111111111100000000000000000000;
11'd1925: out <= 32'b00110000000011000011000000001100;
11'd1926: out <= 32'b00110000000011000011111111110000;
11'd1927: out <= 32'b00000000000000000011111111110000;
11'd1928: out <= 32'b00000011111100000000000000000000;
11'd1929: out <= 32'b00110000000000000000110000001100;
11'd1930: out <= 32'b00001100000011000011000000000000;
11'd1931: out <= 32'b00000000000000000000001111110000;
11'd1932: out <= 32'b00111111110000000000000000000000;
11'd1933: out <= 32'b00110000000011000011000000110000;
11'd1934: out <= 32'b00110000001100000011000000001100;
11'd1935: out <= 32'b00000000000000000011111111000000;
11'd1936: out <= 32'b00111111111111000000000000000000;
11'd1937: out <= 32'b00110000000000000011000000000000;
11'd1938: out <= 32'b00110000000000000011111111000000;
11'd1939: out <= 32'b00000000000000000011000000000000;
11'd1940: out <= 32'b00000011111111000000000000000000;
11'd1941: out <= 32'b00110000000000000000110000000000;
11'd1942: out <= 32'b00001100000011000011000000111100;
11'd1943: out <= 32'b00000000000000000000001111110000;
11'd1944: out <= 32'b00110000000011000000000000000000;
11'd1945: out <= 32'b00110000000011000011000000001100;
11'd1946: out <= 32'b00110000000011000011111111111100;
11'd1947: out <= 32'b00000000000000000011000000001100;
11'd1948: out <= 32'b00000011111100000000000000000000;
11'd1949: out <= 32'b00000000110000000000000011000000;
11'd1950: out <= 32'b00000000110000000000000011000000;
11'd1951: out <= 32'b00000000000000000000001111110000;
11'd1952: out <= 32'b00111111111100000000000000000000;
11'd1953: out <= 32'b00000000110000000000000011000000;
11'd1954: out <= 32'b00110000110000000000000011000000;
11'd1955: out <= 32'b00000000000000000000111100000000;
11'd1956: out <= 32'b00111111111100000000000000000000;
11'd1957: out <= 32'b00000000110000000000000011000000;
11'd1958: out <= 32'b00110000110000000000000011000000;
11'd1959: out <= 32'b00000000000000000000111100000000;
11'd1960: out <= 32'b00110000111100000000000000000000;
11'd1961: out <= 32'b00111100000000000011001100000000;
11'd1962: out <= 32'b00110000110000000011001100000000;
11'd1963: out <= 32'b00000000000000000011000000110000;
11'd1964: out <= 32'b00110000000000000000000000000000;
11'd1965: out <= 32'b00110000000000000011000000000000;
11'd1966: out <= 32'b00110000000000000011000000000000;
11'd1967: out <= 32'b00000000000000000011111111110000;
11'd1968: out <= 32'b00001100111100000000000000000000;
11'd1969: out <= 32'b00110011000011000011001100001100;
11'd1970: out <= 32'b00110000000011000011001100001100;
11'd1971: out <= 32'b00000000000000000011000000001100;
11'd1972: out <= 32'b00110000000011000000000000000000;
11'd1973: out <= 32'b00110011000011000011110000001100;
11'd1974: out <= 32'b00110000001111000011000011001100;
11'd1975: out <= 32'b00000000000000000011000000001100;
11'd1976: out <= 32'b00001111111100000000000000000000;
11'd1977: out <= 32'b00110000000011000011000000001100;
11'd1978: out <= 32'b00110000000011000011000000001100;
11'd1979: out <= 32'b00000000000000000000111111110000;
11'd1980: out <= 32'b00111111111100000000000000000000;
11'd1981: out <= 32'b00110000000011000011000000001100;
11'd1982: out <= 32'b00110000000000000011111111110000;
11'd1983: out <= 32'b00000000000000000011000000000000;
11'd1984: out <= 32'b00001111111100000000000000000000;
11'd1985: out <= 32'b00110000000011000011000000001100;
11'd1986: out <= 32'b00110000110011000011000000001100;
11'd1987: out <= 32'b00000000000011000000111111110000;
11'd1988: out <= 32'b00111111110000000000000000000000;
11'd1989: out <= 32'b00110000110000000011000000110000;
11'd1990: out <= 32'b00110000110000000011111100000000;
11'd1991: out <= 32'b00000000000000000011000000110000;
11'd1992: out <= 32'b00001111110000000000000000000000;
11'd1993: out <= 32'b00110000000000000011000000000000;
11'd1994: out <= 32'b00000000001100000000111111000000;
11'd1995: out <= 32'b00000000000000000000111111000000;
11'd1996: out <= 32'b00111111111111000000000000000000;
11'd1997: out <= 32'b00000011000000000000001100000000;
11'd1998: out <= 32'b00000011000000000000001100000000;
11'd1999: out <= 32'b00000000000000000000001100000000;
11'd2000: out <= 32'b00110000000011000000000000000000;
11'd2001: out <= 32'b00110000000011000011000000001100;
11'd2002: out <= 32'b00110000000011000011000000001100;
11'd2003: out <= 32'b00000000000000000000111111110000;
11'd2004: out <= 32'b00110000000011000000000000000000;
11'd2005: out <= 32'b00110000001100000011000000001100;
11'd2006: out <= 32'b00001100001100000000110000110000;
11'd2007: out <= 32'b00000000000000000000001111000000;
11'd2008: out <= 32'b00110000000011000000000000000000;
11'd2009: out <= 32'b00110000110011000011000000001100;
11'd2010: out <= 32'b00110000110011000011000011001100;
11'd2011: out <= 32'b00000000000000000000111100110000;
11'd2012: out <= 32'b00110000000011000000000000000000;
11'd2013: out <= 32'b00001100001100000011000000001100;
11'd2014: out <= 32'b00001100001100000000001111000000;
11'd2015: out <= 32'b00000000000000000011000000001100;
11'd2016: out <= 32'b00110000000011000000000000000000;
11'd2017: out <= 32'b00001100001100000011000000001100;
11'd2018: out <= 32'b00000011110000000000001111000000;
11'd2019: out <= 32'b00000000000000000000001111000000;
11'd2020: out <= 32'b00111111111111000000000000000000;
11'd2021: out <= 32'b00000000001100000000000000001100;
11'd2022: out <= 32'b00000011000000000000000011000000;
11'd2023: out <= 32'b00000000000000000011111111111100;
11'd2024: out <= 32'b00000000000000000000000000000000;
11'd2025: out <= 32'b00000000000000000000000000000000;
11'd2026: out <= 32'b00000000000000000000000000000000;
11'd2027: out <= 32'b00000000000000000000000110000000;
11'd2028: out <= 32'b00000000000000000000000000000000;
11'd2029: out <= 32'b00000000000000000000000000000000;
11'd2030: out <= 32'b00000000000000000000000000000000;
11'd2031: out <= 32'b00000000011000000000000110000000;
11'd2032: out <= 32'b00000000000000000000000000000000;
11'd2033: out <= 32'b00000000000000000000000110000000;
11'd2034: out <= 32'b00000000000000000000000000000000;
11'd2035: out <= 32'b00000000000000000000000110000000;
11'd2036: out <= 32'b00000000000000000000000000000000;
11'd2037: out <= 32'b00000000000000000000000110000000;
11'd2038: out <= 32'b00000000000000000000000000000000;
11'd2039: out <= 32'b00000000011000000000000110000000;
11'd2040: out <= 32'b00001111111100000000000000000000;
11'd2041: out <= 32'b00111111111100000011110000000000;
11'd2042: out <= 32'b00111111111100000011110000000000;
11'd2043: out <= 32'b00000000000000000011000000000000;
11'd2044: out <= 32'b01000110110101111100111010010000;
11'd2045: out <= 32'b01110110111001100110110011011000;
11'd2046: out <= 32'b00111001000111011111001000001001;
11'd2047: out <= 32'b00001100111010110010011110100111;
default: out <= 0;
endcase
endmodule
